//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT69), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT68), .Z(new_n212));
  OAI21_X1  g0012(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT70), .Z(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  INV_X1    g0017(.A(new_n205), .ZN(new_n218));
  INV_X1    g0018(.A(G13), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(KEYINPUT64), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n205), .B2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT66), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n229), .A2(G1), .A3(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n226), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n216), .A2(new_n217), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G226), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT72), .ZN(new_n250));
  INV_X1    g0050(.A(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT71), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G68), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  NOR2_X1   g0057(.A1(new_n232), .A2(G1), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT76), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n230), .A2(new_n228), .B1(new_n218), .B2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n219), .A2(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G150), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n232), .A2(G33), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n267), .B1(new_n201), .B2(new_n232), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n231), .B1(new_n271), .B2(new_n205), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  INV_X1    g0073(.A(new_n262), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n270), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n265), .A2(KEYINPUT78), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT78), .B1(new_n265), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT9), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n278), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT9), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(new_n276), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT73), .B1(new_n288), .B2(new_n227), .ZN(new_n289));
  AND2_X1   g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT73), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n287), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G226), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G274), .A3(new_n287), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT74), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT75), .ZN(new_n299));
  AND2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n271), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(KEYINPUT75), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n202), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n228), .A2(new_n230), .A3(new_n292), .ZN(new_n309));
  INV_X1    g0109(.A(new_n307), .ZN(new_n310));
  INV_X1    g0110(.A(G223), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G222), .B2(new_n312), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n298), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n295), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n284), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n316), .A2(new_n317), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(G190), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n283), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n283), .B2(new_n320), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G226), .A2(G1698), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n241), .B2(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n302), .A2(new_n326), .A3(new_n306), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n309), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(new_n287), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n288), .A2(KEYINPUT73), .A3(new_n227), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n335));
  OAI211_X1 g0135(.A(G238), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n297), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n297), .A2(new_n336), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n309), .B1(new_n327), .B2(new_n328), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT13), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G169), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n337), .A2(new_n340), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(KEYINPUT14), .B1(new_n343), .B2(G179), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n341), .A2(new_n345), .A3(G169), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(KEYINPUT79), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT79), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n337), .B2(new_n340), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n344), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  INV_X1    g0154(.A(new_n266), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n354), .B1(new_n269), .B2(new_n202), .C1(new_n355), .C2(new_n273), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n356), .A2(new_n272), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(KEYINPUT11), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(KEYINPUT11), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT12), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n360), .A2(new_n219), .A3(G1), .ZN(new_n361));
  INV_X1    g0161(.A(new_n354), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n360), .A2(new_n262), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n353), .B1(new_n263), .B2(KEYINPUT12), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n352), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n343), .A2(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n341), .A2(G200), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n241), .A2(G1698), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G238), .B2(G1698), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n309), .B1(new_n310), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G107), .B2(new_n310), .ZN(new_n376));
  INV_X1    g0176(.A(G274), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n289), .B2(new_n293), .ZN(new_n378));
  AOI22_X1  g0178(.A1(G244), .A2(new_n294), .B1(new_n378), .B2(new_n287), .ZN(new_n379));
  AOI21_X1  g0179(.A(G169), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n264), .A2(G77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G20), .A2(G77), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n382), .B1(new_n268), .B2(new_n355), .C1(new_n269), .C2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n272), .B1(new_n202), .B2(new_n274), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n380), .B2(new_n386), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n376), .A2(new_n379), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(G190), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n386), .C1(new_n284), .C2(new_n391), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n319), .A2(new_n392), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n265), .A2(new_n275), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(G169), .C2(new_n319), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n324), .A2(new_n372), .A3(new_n397), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n268), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n262), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n264), .B2(new_n403), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n304), .A2(new_n232), .A3(new_n305), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT80), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n304), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n305), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT81), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n353), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G58), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n353), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n266), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n272), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n307), .B2(new_n232), .ZN(new_n426));
  INV_X1    g0226(.A(new_n412), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n421), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT16), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n425), .A2(new_n430), .A3(KEYINPUT82), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n406), .A2(new_n408), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n412), .B(KEYINPUT81), .ZN(new_n437));
  OAI21_X1  g0237(.A(G68), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n260), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n300), .A2(new_n301), .A3(new_n299), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT75), .B1(new_n304), .B2(new_n305), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n232), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n427), .B1(new_n442), .B2(new_n408), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n429), .B1(new_n443), .B2(new_n353), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n422), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n432), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n405), .B1(new_n431), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n405), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT82), .B1(new_n425), .B2(new_n430), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n439), .A2(new_n445), .A3(new_n432), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n311), .A2(new_n312), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(G226), .B2(new_n312), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n300), .A2(new_n301), .ZN(new_n457));
  INV_X1    g0257(.A(G87), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n456), .A2(new_n457), .B1(new_n271), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n330), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n294), .A2(G232), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n297), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n349), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n392), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n449), .A2(new_n454), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT18), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n449), .A2(new_n470), .A3(new_n454), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(G200), .ZN(new_n472));
  INV_X1    g0272(.A(G190), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n453), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n450), .B(new_n474), .C1(new_n451), .C2(new_n452), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT17), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n469), .A2(new_n471), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n402), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n286), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n296), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(G257), .B1(new_n378), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n302), .A2(new_n306), .A3(G250), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n312), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g0292(.A(G244), .B1(new_n300), .B2(new_n301), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n493), .A2(new_n494), .B1(G33), .B2(G283), .ZN(new_n495));
  INV_X1    g0295(.A(G244), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n494), .A2(new_n496), .A3(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n302), .A2(new_n306), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT84), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n330), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT84), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n490), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT85), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR3_X1    g0305(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT84), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n330), .A3(new_n500), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n490), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n508), .A3(G200), .ZN(new_n509));
  OAI211_X1 g0309(.A(G190), .B(new_n490), .C1(new_n501), .C2(new_n502), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n274), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G1), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G33), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n260), .A2(new_n262), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n515), .B2(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n248), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n511), .A2(new_n248), .ZN(new_n518));
  NOR2_X1   g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(KEYINPUT6), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n443), .B2(new_n248), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n516), .B1(new_n523), .B2(new_n272), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n507), .A2(new_n392), .A3(new_n490), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n503), .B2(new_n349), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n509), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(G250), .B1(new_n513), .B2(G45), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n377), .B2(new_n485), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n296), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G238), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n496), .B2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n304), .A2(new_n305), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G33), .B2(G116), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n531), .B(G190), .C1(new_n535), .C2(new_n309), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n309), .ZN(new_n537));
  INV_X1    g0337(.A(new_n531), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(new_n284), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n458), .A2(new_n511), .A3(new_n248), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n328), .A2(new_n232), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT19), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n232), .B(G68), .C1(new_n300), .C2(new_n301), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n269), .B2(new_n511), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT86), .A4(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n272), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n274), .A2(new_n383), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n458), .C2(new_n515), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n540), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n515), .ZN(new_n555));
  INV_X1    g0355(.A(new_n383), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n557), .A3(new_n552), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n260), .B1(new_n547), .B2(new_n548), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n550), .B1(new_n274), .B2(new_n383), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(KEYINPUT87), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n535), .A2(new_n309), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(G179), .A3(new_n531), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n539), .B2(new_n349), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n554), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n458), .A2(KEYINPUT22), .A3(G20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n302), .A2(new_n306), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT89), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT89), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n534), .A2(new_n232), .A3(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n248), .A2(KEYINPUT23), .A3(G20), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT23), .B1(new_n248), .B2(G20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G116), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n580), .A2(new_n581), .B1(G20), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n569), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n573), .A2(new_n574), .B1(KEYINPUT22), .B2(new_n576), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(KEYINPUT24), .A3(new_n583), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n272), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n274), .B(new_n248), .C1(KEYINPUT90), .C2(KEYINPUT25), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n555), .A2(G107), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G257), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G1698), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G250), .B2(G1698), .ZN(new_n597));
  INV_X1    g0397(.A(G294), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n597), .A2(new_n457), .B1(new_n271), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n330), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n378), .A2(new_n489), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n296), .A2(G264), .A3(new_n487), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n473), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT91), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n284), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(KEYINPUT91), .A3(new_n284), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n588), .A2(new_n594), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n568), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n528), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n260), .A2(G116), .A3(new_n262), .A4(new_n514), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n274), .A2(new_n251), .ZN(new_n614));
  AOI21_X1  g0414(.A(G20), .B1(G33), .B2(G283), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n271), .A2(G97), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(G20), .B2(new_n251), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT20), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n260), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n272), .B2(new_n617), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n613), .B(new_n614), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT88), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G264), .A2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n457), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n534), .A2(KEYINPUT88), .A3(G264), .A4(G1698), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n534), .A2(G257), .A3(new_n312), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G303), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n302), .B2(new_n306), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n330), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n488), .A2(G270), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n601), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n622), .B1(new_n633), .B2(G200), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n473), .B2(new_n633), .ZN(new_n635));
  INV_X1    g0435(.A(new_n633), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(G179), .A3(new_n622), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n622), .A2(G169), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT21), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n619), .B1(new_n618), .B2(new_n260), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n272), .A2(KEYINPUT20), .A3(new_n617), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n251), .B2(new_n274), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n349), .B1(new_n643), .B2(new_n613), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n644), .B2(new_n633), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n635), .B(new_n637), .C1(new_n639), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n605), .A2(G179), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n605), .A2(new_n349), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n578), .A2(new_n569), .A3(new_n584), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT24), .B1(new_n586), .B2(new_n583), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n260), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n647), .B(new_n648), .C1(new_n651), .C2(new_n593), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n483), .A2(new_n612), .A3(new_n654), .ZN(G372));
  OAI21_X1  g0455(.A(new_n637), .B1(new_n639), .B2(new_n645), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT92), .ZN(new_n657));
  INV_X1    g0457(.A(new_n622), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n658), .A2(new_n633), .A3(new_n392), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT21), .B1(new_n636), .B2(new_n638), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n644), .A2(new_n640), .A3(new_n633), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n657), .A2(new_n664), .A3(new_n652), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n528), .A3(new_n611), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n558), .A2(new_n559), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT87), .B1(new_n562), .B2(new_n557), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n567), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n503), .A2(new_n349), .ZN(new_n672));
  INV_X1    g0472(.A(new_n524), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n526), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n554), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n568), .A2(KEYINPUT26), .A3(new_n526), .A4(new_n527), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n670), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n666), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n483), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n447), .A2(new_n470), .A3(new_n467), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT18), .B1(new_n453), .B2(new_n466), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n371), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n394), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n367), .B2(new_n352), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n453), .A2(new_n479), .A3(new_n475), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n479), .B1(new_n453), .B2(new_n475), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n685), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n324), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n401), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n681), .A2(new_n694), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n261), .A2(new_n232), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(G213), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n588), .B2(new_n594), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT94), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n610), .A3(new_n652), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(KEYINPUT94), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n653), .B2(new_n701), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n657), .A2(new_n664), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n658), .A2(new_n702), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n646), .B(KEYINPUT93), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(G330), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT95), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n662), .A2(new_n701), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n653), .A2(new_n702), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n716), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n223), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n541), .A2(G116), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n723), .A2(new_n513), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n235), .B2(new_n723), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT28), .Z(new_n727));
  NAND2_X1  g0527(.A1(new_n680), .A2(new_n702), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n662), .A2(new_n652), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n509), .A2(new_n525), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n611), .A2(new_n730), .A3(new_n731), .A4(new_n674), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n701), .B1(new_n679), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n631), .A2(new_n632), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n566), .A2(new_n605), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n507), .A2(new_n490), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n539), .A2(G179), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n742), .A2(new_n633), .A3(new_n605), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(new_n741), .B1(new_n503), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n738), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n745), .A2(new_n503), .A3(new_n741), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n702), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(new_n747), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n654), .A2(new_n528), .A3(new_n611), .A4(new_n702), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n737), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n736), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n727), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n714), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n219), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n513), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n723), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n722), .A2(new_n307), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n768), .A2(G355), .B1(new_n251), .B2(new_n722), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n256), .A2(G45), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n722), .A2(new_n534), .ZN(new_n771));
  INV_X1    g0571(.A(new_n235), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(G45), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n231), .B1(G20), .B2(new_n349), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n760), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n767), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n232), .A2(G179), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(G329), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n232), .A2(new_n392), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G190), .A3(new_n284), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n473), .A2(new_n284), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(G322), .B1(new_n791), .B2(G326), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n473), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n232), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n307), .C1(new_n598), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n789), .A2(new_n778), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n284), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n778), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n796), .A2(new_n629), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  NAND2_X1  g0601(.A1(new_n786), .A2(new_n797), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n786), .A2(new_n779), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n785), .A2(new_n795), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n796), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G87), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n310), .B(new_n808), .C1(new_n248), .C2(new_n798), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT99), .ZN(new_n810));
  INV_X1    g0610(.A(new_n803), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n202), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n794), .A2(new_n511), .ZN(new_n817));
  INV_X1    g0617(.A(new_n802), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G50), .A2(new_n791), .B1(new_n818), .B2(G68), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n416), .B2(new_n787), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n810), .A2(new_n816), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n783), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT32), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n806), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n775), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n777), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n762), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n714), .A2(G330), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n714), .A2(G330), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n767), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n386), .A2(new_n702), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n394), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n394), .A2(KEYINPUT103), .A3(new_n396), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n394), .A2(new_n838), .A3(new_n396), .ZN(new_n839));
  INV_X1    g0639(.A(new_n835), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n836), .A2(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n728), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n701), .B1(new_n666), .B2(new_n679), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n753), .A3(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT104), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n767), .B1(new_n753), .B2(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n798), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n457), .B1(new_n852), .B2(G68), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n273), .B2(new_n796), .C1(new_n416), .C2(new_n794), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n788), .A2(G143), .B1(new_n818), .B2(G150), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n856), .B2(new_n790), .C1(new_n815), .C2(new_n822), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  AOI211_X1 g0658(.A(new_n854), .B(new_n858), .C1(G132), .C2(new_n784), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n787), .A2(new_n598), .B1(new_n802), .B2(new_n799), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n790), .A2(new_n629), .B1(new_n796), .B2(new_n248), .ZN(new_n861));
  OR4_X1    g0661(.A1(new_n310), .A2(new_n860), .A3(new_n861), .A4(new_n817), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(G87), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n783), .B2(new_n804), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT102), .ZN(new_n865));
  INV_X1    g0665(.A(new_n815), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n862), .B(new_n865), .C1(G116), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n775), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n775), .A2(new_n758), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n767), .B1(new_n869), .B2(new_n202), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n868), .B(new_n870), .C1(new_n841), .C2(new_n759), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n851), .A2(new_n871), .ZN(G384));
  NOR2_X1   g0672(.A1(new_n763), .A2(new_n513), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n749), .B1(new_n747), .B2(KEYINPUT110), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT110), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n876), .B(new_n702), .C1(new_n744), .C2(new_n746), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n752), .B(new_n874), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n367), .A2(new_n701), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n337), .A2(new_n340), .A3(G179), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n350), .B2(new_n345), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n346), .A2(KEYINPUT79), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n350), .A2(new_n348), .A3(new_n345), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n371), .B(new_n879), .C1(new_n884), .C2(new_n366), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT106), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n368), .A2(new_n887), .A3(new_n371), .A4(new_n879), .ZN(new_n888));
  INV_X1    g0688(.A(new_n879), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n886), .A2(new_n888), .B1(new_n352), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n842), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n438), .B2(new_n429), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n405), .B1(new_n425), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n699), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n893), .A2(KEYINPUT107), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT107), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n468), .A2(KEYINPUT18), .B1(new_n477), .B2(new_n480), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n471), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n453), .A2(new_n475), .B1(new_n467), .B2(new_n893), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n476), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n448), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(new_n467), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n449), .A2(new_n454), .A3(new_n894), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n899), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n469), .A2(new_n471), .A3(new_n481), .ZN(new_n913));
  INV_X1    g0713(.A(new_n897), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n902), .ZN(new_n916));
  INV_X1    g0716(.A(new_n903), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n478), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n468), .A2(new_n909), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n878), .B(new_n891), .C1(new_n912), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n920), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n905), .A2(new_n906), .A3(new_n699), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n691), .B2(new_n684), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n468), .A2(new_n909), .A3(new_n918), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n453), .A2(new_n466), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n478), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n903), .B1(new_n909), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n911), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n352), .A2(new_n889), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n686), .B1(new_n352), .B2(new_n367), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n887), .B1(new_n935), .B2(new_n879), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND4_X1   g0738(.A1(KEYINPUT40), .A2(new_n938), .A3(new_n878), .A4(new_n841), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n922), .A2(new_n923), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n483), .A2(new_n878), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n737), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT111), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n368), .A2(new_n701), .ZN(new_n946));
  XNOR2_X1  g0746(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n924), .A2(new_n932), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n911), .B1(new_n899), .B2(new_n910), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n924), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n685), .A2(new_n894), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n924), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n394), .A2(new_n701), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n844), .B2(new_n841), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n890), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n483), .B1(new_n729), .B2(new_n735), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n694), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n873), .B1(new_n945), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n945), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n965));
  OAI211_X1 g0765(.A(G116), .B(new_n233), .C1(new_n521), .C2(KEYINPUT35), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT105), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT36), .Z(new_n970));
  NOR3_X1   g0770(.A1(new_n772), .A2(new_n202), .A3(new_n417), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n353), .A2(G50), .ZN(new_n972));
  OAI211_X1 g0772(.A(G1), .B(new_n219), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n964), .A2(new_n970), .A3(new_n973), .ZN(G367));
  OAI21_X1  g0774(.A(new_n528), .B1(new_n524), .B2(new_n702), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n527), .A2(new_n526), .A3(new_n701), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n707), .A3(new_n717), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n674), .B1(new_n975), .B2(new_n652), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n978), .A2(KEYINPUT42), .B1(new_n702), .B2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n553), .A2(new_n701), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n676), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n670), .A2(new_n982), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n979), .A2(new_n981), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n988), .B(new_n989), .Z(new_n990));
  INV_X1    g0790(.A(new_n716), .ZN(new_n991));
  INV_X1    g0791(.A(new_n977), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n990), .B(new_n993), .Z(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n723), .B(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n720), .A2(new_n992), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n720), .A2(new_n992), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT44), .Z(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n998), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n716), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n718), .B1(new_n709), .B2(new_n717), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n831), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n755), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n996), .B1(new_n1010), .B2(new_n756), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n994), .B1(new_n1011), .B2(new_n765), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n771), .A2(new_n245), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n776), .B1(new_n223), .B2(new_n383), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n766), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G294), .A2(new_n818), .B1(new_n852), .B2(G97), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n629), .B2(new_n787), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n815), .A2(new_n799), .B1(new_n1018), .B2(new_n783), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n457), .B1(new_n790), .B2(new_n804), .C1(new_n794), .C2(new_n248), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT114), .B1(new_n796), .B2(new_n251), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT46), .ZN(new_n1022));
  OR4_X1    g0822(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G58), .A2(new_n807), .B1(new_n818), .B2(G159), .ZN(new_n1024));
  INV_X1    g0824(.A(G150), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n787), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n866), .B2(G50), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n852), .A2(G77), .ZN(new_n1028));
  INV_X1    g0828(.A(G143), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n790), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n794), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n307), .B(new_n1030), .C1(G68), .C2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1027), .B(new_n1032), .C1(new_n856), .C2(new_n783), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1023), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n775), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n987), .B2(new_n761), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT115), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n1012), .A2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n1009), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1008), .A2(new_n755), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n723), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n202), .A2(new_n796), .B1(new_n802), .B2(new_n268), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n457), .B(new_n1043), .C1(G97), .C2(new_n852), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1031), .A2(new_n556), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n784), .A2(G150), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n787), .A2(new_n273), .B1(new_n790), .B2(new_n822), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G68), .B2(new_n811), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n784), .A2(G326), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n534), .B1(new_n852), .B2(G116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n794), .A2(new_n799), .B1(new_n796), .B2(new_n598), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G322), .A2(new_n791), .B1(new_n818), .B2(G311), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n1018), .B2(new_n787), .C1(new_n815), .C2(new_n629), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1050), .B(new_n1051), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n775), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n242), .A2(G45), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1063), .A2(new_n771), .B1(new_n724), .B2(new_n768), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n403), .A2(new_n273), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n286), .B1(new_n353), .B2(new_n202), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1066), .A2(new_n724), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1064), .A2(new_n1068), .B1(G107), .B2(new_n223), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n767), .B1(new_n1069), .B2(new_n776), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1062), .B(new_n1070), .C1(new_n709), .C2(new_n761), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1042), .B(new_n1071), .C1(new_n764), .C2(new_n1008), .ZN(G393));
  OAI21_X1  g0872(.A(new_n1040), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1010), .A2(new_n723), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n992), .A2(new_n760), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n815), .A2(new_n268), .B1(new_n273), .B2(new_n802), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT116), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n787), .A2(new_n822), .B1(new_n790), .B2(new_n1025), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1031), .A2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n807), .A2(G68), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1080), .A2(new_n534), .A3(new_n863), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G143), .B2(new_n784), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1077), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n787), .A2(new_n804), .B1(new_n790), .B2(new_n1018), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n784), .A2(G322), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n799), .A2(new_n796), .B1(new_n802), .B2(new_n629), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n803), .A2(new_n598), .B1(new_n798), .B2(new_n248), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n310), .B1(G116), .B2(new_n1031), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n826), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n776), .B1(new_n511), .B2(new_n223), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n252), .B2(new_n771), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n767), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1006), .A2(new_n765), .B1(new_n1075), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1074), .A2(new_n1097), .ZN(G390));
  OAI21_X1  g0898(.A(KEYINPUT39), .B1(new_n912), .B2(new_n921), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n924), .A2(new_n932), .A3(new_n947), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n946), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n956), .B2(new_n890), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n753), .A2(new_n841), .A3(new_n938), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n955), .B1(new_n733), .B2(new_n841), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n933), .B(new_n1101), .C1(new_n890), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n677), .A2(new_n678), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n732), .A2(new_n1108), .A3(new_n669), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n841), .A3(new_n702), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n955), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n890), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n946), .B(new_n1112), .C1(new_n924), .C2(new_n932), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n948), .A2(new_n951), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n1102), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n891), .A2(G330), .A3(new_n878), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n765), .B(new_n1107), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT118), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n948), .A2(new_n951), .A3(new_n759), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n869), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n852), .A2(G68), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1080), .A2(new_n307), .A3(new_n808), .A4(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n788), .A2(G116), .B1(new_n818), .B2(G107), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n799), .B2(new_n790), .C1(new_n815), .C2(new_n511), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(G294), .C2(new_n784), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n310), .B1(new_n273), .B2(new_n798), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n784), .B2(G125), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n1025), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT53), .B1(new_n796), .B2(new_n1025), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n822), .C2(new_n794), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n788), .A2(G132), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1132), .B1(new_n802), .B2(new_n856), .C1(new_n1133), .C2(new_n790), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1131), .B(new_n1134), .C1(new_n866), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1125), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n766), .B1(new_n403), .B2(new_n1120), .C1(new_n1138), .C2(new_n826), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1119), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1117), .A2(new_n1118), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1118), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1116), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n764), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT118), .B1(new_n1147), .B2(new_n1140), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1117), .A2(new_n1118), .A3(new_n1141), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n956), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1116), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n938), .B1(new_n753), .B2(new_n841), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n878), .A2(G330), .A3(new_n841), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1104), .B(new_n1105), .C1(new_n1156), .C2(new_n938), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n483), .A2(G330), .A3(new_n878), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n960), .A2(new_n1159), .A3(new_n694), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1107), .B(new_n1164), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1165), .A3(new_n723), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1144), .A2(new_n1151), .A3(new_n1166), .ZN(G378));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n693), .B2(new_n400), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n699), .B1(new_n280), .B2(new_n276), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n324), .A2(new_n401), .A3(new_n1168), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n940), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n909), .A2(new_n929), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n919), .B1(new_n1178), .B2(new_n903), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT38), .B1(new_n1179), .B2(new_n926), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n939), .B1(new_n912), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n938), .A2(new_n878), .A3(new_n841), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n950), .B2(new_n924), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(G330), .C1(new_n1183), .C2(KEYINPUT40), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT123), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n959), .B2(KEYINPUT122), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT122), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1189), .B(KEYINPUT123), .C1(new_n952), .C2(new_n958), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1186), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1184), .B(new_n1176), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1101), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n954), .A2(new_n957), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n953), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT122), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT123), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n959), .A2(KEYINPUT122), .A3(new_n1187), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1192), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1165), .A2(new_n1161), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1191), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n723), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1186), .A2(new_n959), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1177), .A2(new_n952), .A3(new_n1185), .A4(new_n958), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1203), .B1(new_n1165), .B2(new_n1161), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1205), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1204), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1191), .A2(new_n1200), .A3(new_n765), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n285), .B(new_n457), .C1(new_n796), .C2(new_n202), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n787), .A2(new_n248), .B1(new_n790), .B2(new_n251), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G68), .C2(new_n1031), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n803), .A2(new_n383), .B1(new_n798), .B2(new_n416), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G97), .B2(new_n818), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(new_n799), .C2(new_n783), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT58), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n273), .B1(new_n300), .B2(G41), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n787), .A2(new_n1133), .B1(new_n803), .B2(new_n856), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G125), .B2(new_n791), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G132), .A2(new_n818), .B1(new_n807), .B2(new_n1136), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n1025), .C2(new_n794), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n784), .A2(G124), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G33), .B(G41), .C1(new_n852), .C2(G159), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1219), .B(new_n1220), .C1(new_n1225), .C2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n775), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT121), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n767), .B1(new_n869), .B2(new_n273), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n1176), .C2(new_n759), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1212), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1211), .A2(new_n1236), .ZN(G375));
  NAND3_X1  g1037(.A1(new_n1155), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n996), .B(KEYINPUT124), .Z(new_n1239));
  NAND3_X1  g1039(.A1(new_n1162), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n890), .A2(new_n758), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n766), .B1(G68), .B2(new_n1120), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n790), .A2(new_n598), .B1(new_n796), .B2(new_n511), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G116), .B2(new_n818), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n629), .B2(new_n783), .C1(new_n815), .C2(new_n248), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n788), .A2(G283), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1045), .A2(new_n1246), .A3(new_n307), .A4(new_n1028), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G150), .A2(new_n811), .B1(new_n807), .B2(G159), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n457), .B1(new_n852), .B2(G58), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n273), .C2(new_n794), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n788), .A2(G137), .B1(new_n791), .B2(G132), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n802), .B2(new_n1135), .C1(new_n1133), .C2(new_n783), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1245), .A2(new_n1247), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1242), .B1(new_n1253), .B2(new_n775), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1158), .A2(new_n765), .B1(new_n1241), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1240), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1012), .A3(new_n1038), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G381), .ZN(new_n1259));
  INV_X1    g1059(.A(G375), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1166), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT125), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .A4(new_n1265), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n700), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1260), .A2(new_n1263), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  NAND2_X1  g1070(.A1(G387), .A2(G390), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(G396), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1271), .A2(new_n1258), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1271), .B2(new_n1258), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G378), .A2(new_n1211), .A3(new_n1236), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1208), .A2(new_n765), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1239), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1279), .B(new_n1235), .C1(new_n1202), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1263), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1238), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1155), .A2(new_n1160), .A3(KEYINPUT60), .A4(new_n1157), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n723), .A3(new_n1162), .A4(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G384), .A3(new_n1255), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1287), .B2(new_n1255), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1283), .A2(new_n1267), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1276), .B1(new_n1277), .B2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1277), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1268), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G2897), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1267), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1300), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1303), .B2(new_n1298), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1295), .B1(new_n1296), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1294), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1293), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1292), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1296), .A2(KEYINPUT62), .A3(new_n1291), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1305), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1276), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1283), .A2(new_n1267), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1303), .A2(new_n1298), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1291), .A2(new_n1297), .A3(new_n1302), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1310), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT62), .B1(new_n1296), .B2(new_n1291), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1318), .B(new_n1312), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1307), .B1(new_n1313), .B2(new_n1322), .ZN(G405));
  INV_X1    g1123(.A(new_n1263), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1278), .B1(new_n1260), .B2(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1291), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1276), .ZN(G402));
endmodule


