//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n188), .A2(new_n190), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  INV_X1    g014(.A(G110), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G128), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  XNOR2_X1  g018(.A(G119), .B(G128), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n203), .A2(KEYINPUT73), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n193), .B(new_n195), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(new_n202), .A3(new_n200), .ZN(new_n209));
  AOI22_X1  g023(.A1(G110), .A2(new_n209), .B1(new_n204), .B2(new_n205), .ZN(new_n210));
  INV_X1    g024(.A(new_n193), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G137), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n215), .A2(KEYINPUT74), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(KEYINPUT74), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  OR3_X1    g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n216), .B2(new_n217), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n208), .A3(new_n213), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n229), .A3(new_n224), .A4(new_n226), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(G234), .B2(new_n224), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT75), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n228), .A2(new_n235), .A3(new_n230), .A4(new_n232), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(G902), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G472), .ZN(new_n240));
  NOR2_X1   g054(.A1(G237), .A2(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G210), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n242), .B(KEYINPUT27), .Z(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT71), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT26), .B(G101), .Z(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT11), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n254), .A2(new_n255), .A3(new_n257), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n257), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT66), .A3(G131), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  XNOR2_X1  g079(.A(G134), .B(G137), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n255), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT1), .B1(new_n269), .B2(G146), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(G146), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n194), .A2(G143), .ZN(new_n272));
  OAI211_X1 g086(.A(G128), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n194), .A2(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(G146), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(new_n275), .C1(KEYINPUT1), .C2(new_n199), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n260), .B1(new_n258), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n257), .B1(new_n253), .B2(new_n250), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  XNOR2_X1  g097(.A(G143), .B(G146), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT0), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n199), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT0), .B(G128), .Z(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n267), .A2(new_n264), .ZN(new_n290));
  INV_X1    g104(.A(new_n277), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n262), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n278), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  INV_X1    g109(.A(G116), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(G119), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n197), .A2(G116), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT2), .B(G113), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n197), .A2(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(G119), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT2), .B(G113), .Z(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(KEYINPUT70), .A3(new_n301), .A4(new_n302), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n302), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n300), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n299), .A2(KEYINPUT69), .A3(new_n300), .A4(new_n303), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n294), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n262), .A2(new_n264), .A3(new_n267), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n316), .A2(new_n291), .B1(new_n283), .B2(new_n288), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n306), .A2(new_n313), .A3(new_n312), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n248), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n248), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n247), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n324));
  NAND2_X1  g138(.A1(new_n294), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(KEYINPUT30), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n314), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n246), .A4(new_n319), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n268), .A2(new_n277), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n287), .A2(new_n284), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n282), .A2(new_n262), .B1(new_n332), .B2(new_n286), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n331), .A2(new_n314), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n294), .A2(new_n324), .B1(new_n317), .B2(KEYINPUT30), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n314), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n328), .B1(new_n336), .B2(new_n246), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n240), .B(new_n224), .C1(new_n330), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT32), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n327), .A2(new_n246), .A3(new_n319), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT31), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n329), .A3(new_n323), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n240), .A4(new_n224), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n334), .B1(new_n314), .B2(new_n294), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n246), .B(new_n321), .C1(new_n347), .C2(new_n248), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n336), .A2(new_n246), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n327), .A2(new_n319), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n247), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n349), .A4(new_n348), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n317), .B(new_n318), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n322), .B1(new_n356), .B2(KEYINPUT28), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n247), .A2(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G472), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n239), .B1(new_n345), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT9), .B(G234), .ZN(new_n363));
  OAI21_X1  g177(.A(G221), .B1(new_n363), .B2(G902), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT76), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n369), .A2(G104), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n371), .A2(new_n372), .A3(new_n374), .A4(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n373), .B2(new_n376), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT78), .B1(new_n382), .B2(new_n277), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT10), .ZN(new_n384));
  INV_X1    g198(.A(new_n283), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT78), .B(new_n386), .C1(new_n382), .C2(new_n277), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n371), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n372), .B1(new_n388), .B2(new_n371), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n288), .B(new_n391), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n384), .A2(new_n385), .A3(new_n387), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n282), .B2(new_n262), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n382), .A2(new_n277), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n380), .A2(new_n381), .B1(new_n276), .B2(new_n273), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT12), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT12), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n395), .A2(new_n401), .A3(KEYINPUT80), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n218), .A2(G227), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n401), .A3(new_n403), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n395), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n387), .A2(new_n394), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n291), .A2(new_n381), .A3(new_n380), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n386), .B1(new_n415), .B2(KEYINPUT78), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n283), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n409), .A2(new_n412), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G469), .B1(new_n418), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n395), .A2(new_n401), .A3(new_n403), .A4(new_n407), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n407), .B1(new_n417), .B2(new_n395), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n420), .B(new_n224), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n395), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n408), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n420), .A4(new_n224), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n365), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  INV_X1    g247(.A(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n218), .A3(G214), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n241), .B(G214), .C1(new_n436), .C2(G143), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n433), .B(new_n255), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n255), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n255), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n443), .B2(new_n433), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n211), .B2(new_n212), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n191), .A2(new_n192), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n194), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT89), .A3(new_n193), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n375), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n438), .A2(new_n439), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT18), .A2(G131), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n194), .B1(new_n188), .B2(new_n190), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n195), .ZN(new_n462));
  INV_X1    g276(.A(new_n195), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(new_n460), .A3(KEYINPUT87), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n457), .B(new_n458), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n453), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(G131), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n438), .A2(new_n439), .A3(new_n255), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT19), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT19), .B1(new_n188), .B2(new_n190), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n194), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n194), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n469), .A2(new_n473), .A3(new_n193), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n465), .ZN(new_n477));
  INV_X1    g291(.A(new_n453), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT90), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n485), .A3(new_n481), .A4(new_n482), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n453), .B1(new_n476), .B2(new_n465), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n462), .A2(new_n464), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n455), .A2(new_n456), .B1(new_n442), .B2(KEYINPUT18), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n444), .A2(new_n450), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n490), .B2(new_n453), .ZN(new_n491));
  INV_X1    g305(.A(new_n482), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT20), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n486), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n451), .A2(new_n465), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n478), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n496), .B2(new_n466), .ZN(new_n497));
  INV_X1    g311(.A(G475), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G128), .B(G143), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n502), .A2(G134), .ZN(new_n503));
  INV_X1    g317(.A(G122), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G116), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n296), .A2(G122), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n369), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(G134), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n510), .B(KEYINPUT14), .C1(new_n504), .C2(G116), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n296), .A3(G122), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n506), .B2(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g329(.A(G107), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT94), .B(G107), .C1(new_n514), .C2(new_n515), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n509), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n199), .A2(G143), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n256), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n502), .ZN(new_n524));
  INV_X1    g338(.A(new_n507), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n369), .B1(new_n505), .B2(new_n506), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n505), .A2(new_n506), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT91), .B1(new_n530), .B2(new_n507), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n524), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n527), .B1(new_n525), .B2(new_n526), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(KEYINPUT91), .A3(new_n507), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n524), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n520), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n363), .A2(new_n231), .A3(G953), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT95), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n518), .A2(new_n519), .ZN(new_n542));
  INV_X1    g356(.A(new_n509), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n524), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT92), .B1(new_n537), .B2(new_n524), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n548));
  INV_X1    g362(.A(new_n540), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n539), .A2(new_n540), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n541), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n224), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n224), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(G234), .A2(G237), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G952), .A3(new_n218), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT96), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n560), .A2(G902), .A3(G953), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n501), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n382), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT5), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n197), .A3(G116), .ZN(new_n570));
  OAI21_X1  g384(.A(G113), .B1(new_n570), .B2(KEYINPUT82), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(KEYINPUT82), .B2(new_n570), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT68), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT68), .B1(new_n301), .B2(new_n302), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT5), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n576), .A3(new_n312), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n318), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G110), .B(G122), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT83), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n577), .B(new_n581), .C1(new_n318), .C2(new_n578), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n586), .A3(new_n582), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n277), .A2(new_n189), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n189), .B2(new_n288), .ZN(new_n589));
  INV_X1    g403(.A(G224), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G953), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n585), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n576), .A2(new_n312), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n581), .A2(KEYINPUT8), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n581), .A2(KEYINPUT8), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n594), .A2(new_n382), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n572), .B1(new_n569), .B2(new_n310), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n312), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n568), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n601));
  OAI221_X1 g415(.A(new_n588), .B1(new_n601), .B2(new_n591), .C1(new_n189), .C2(new_n288), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n589), .B(KEYINPUT7), .C1(new_n590), .C2(G953), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n597), .A2(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n604), .B2(new_n584), .ZN(new_n605));
  OAI21_X1  g419(.A(G210), .B1(G237), .B2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n593), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n593), .A2(new_n605), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n606), .B(KEYINPUT84), .Z(new_n609));
  AOI21_X1  g423(.A(KEYINPUT85), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT85), .ZN(new_n611));
  INV_X1    g425(.A(new_n609), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n611), .B(new_n612), .C1(new_n593), .C2(new_n605), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(G214), .B1(G237), .B2(G902), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n362), .A2(new_n432), .A3(new_n567), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(new_n566), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n593), .A2(new_n605), .A3(new_n606), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n606), .B1(new_n593), .B2(new_n605), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n619), .B(new_n615), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n552), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n547), .B2(new_n549), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n551), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n554), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n553), .A2(new_n554), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n501), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n629), .A2(new_n630), .B1(new_n494), .B2(new_n500), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT98), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n622), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n338), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n240), .B1(new_n342), .B2(new_n224), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n239), .B(new_n365), .C1(new_n419), .C2(new_n431), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  INV_X1    g459(.A(new_n466), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n453), .B1(new_n451), .B2(new_n465), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n224), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n493), .A2(new_n483), .B1(new_n648), .B2(G475), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n559), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n645), .B1(new_n622), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n615), .ZN(new_n652));
  INV_X1    g466(.A(new_n606), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n608), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n654), .B2(new_n607), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n481), .B1(new_n480), .B2(new_n482), .ZN(new_n656));
  AOI211_X1 g470(.A(KEYINPUT20), .B(new_n492), .C1(new_n466), .C2(new_n479), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n656), .A2(new_n657), .B1(new_n497), .B2(new_n498), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n556), .B2(new_n558), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(KEYINPUT99), .A3(new_n659), .A4(new_n619), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n640), .A3(new_n641), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  OAI21_X1  g478(.A(new_n224), .B1(new_n330), .B2(new_n337), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n214), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n237), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n234), .A2(new_n236), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n234), .A2(KEYINPUT100), .A3(new_n236), .A4(new_n669), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n666), .A2(new_n338), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n616), .A3(new_n432), .A4(new_n567), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n563), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT101), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT101), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n562), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n655), .A2(new_n679), .A3(new_n659), .A4(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n552), .A2(new_n224), .A3(new_n557), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n557), .B1(new_n552), .B2(new_n224), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n649), .B(new_n686), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT103), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n687), .A2(new_n692), .A3(new_n432), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n672), .A2(new_n673), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n345), .B2(new_n361), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XOR2_X1   g511(.A(new_n685), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n432), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n614), .A2(KEYINPUT38), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n614), .A2(KEYINPUT38), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n501), .A2(new_n559), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n652), .A3(new_n670), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n340), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n247), .B2(new_n356), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n345), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT104), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n269), .ZN(G45));
  NAND3_X1  g528(.A1(new_n631), .A2(new_n501), .A3(new_n686), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n688), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n695), .A2(new_n432), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  INV_X1    g532(.A(new_n365), .ZN(new_n719));
  INV_X1    g533(.A(new_n428), .ZN(new_n720));
  OAI21_X1  g534(.A(G469), .B1(new_n720), .B2(G902), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n431), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n637), .A2(new_n362), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n362), .A2(new_n661), .A3(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n722), .A2(new_n688), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n695), .A2(new_n567), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  OAI21_X1  g545(.A(new_n329), .B1(new_n357), .B2(new_n246), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n240), .B(new_n224), .C1(new_n732), .C2(new_n337), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n666), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n239), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n705), .A2(new_n688), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n619), .A3(new_n723), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR3_X1   g552(.A1(new_n722), .A2(new_n715), .A3(new_n688), .ZN(new_n739));
  INV_X1    g553(.A(new_n670), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  AND2_X1   g557(.A1(new_n419), .A2(new_n431), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n615), .B(new_n607), .C1(new_n610), .C2(new_n613), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n365), .ZN(new_n746));
  INV_X1    g560(.A(new_n715), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n362), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n746), .A2(new_n362), .A3(KEYINPUT42), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  XNOR2_X1  g567(.A(new_n691), .B(KEYINPUT105), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n746), .A2(new_n362), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND2_X1  g570(.A1(new_n413), .A2(new_n417), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n410), .A2(new_n411), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n404), .A2(new_n408), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  NAND2_X1  g576(.A1(G469), .A2(G902), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n765), .B(G469), .C1(new_n761), .C2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n431), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n719), .A3(new_n698), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n640), .A2(new_n740), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n631), .A2(new_n500), .A3(new_n494), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT43), .ZN(new_n773));
  INV_X1    g587(.A(new_n501), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n631), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n770), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n768), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n777), .A4(new_n773), .ZN(new_n780));
  INV_X1    g594(.A(new_n745), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT107), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT107), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  NAND2_X1  g600(.A1(new_n767), .A2(new_n719), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n719), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n339), .A2(new_n344), .B1(new_n360), .B2(G472), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n792), .A2(new_n239), .A3(new_n747), .A4(new_n781), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n670), .A2(new_n685), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n711), .A2(new_n432), .A3(new_n736), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n696), .A2(new_n717), .A3(new_n742), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n693), .A2(new_n695), .B1(new_n739), .B2(new_n741), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .A3(new_n717), .A4(new_n799), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n724), .A2(new_n727), .A3(new_n730), .A4(new_n737), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  INV_X1    g621(.A(new_n239), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n640), .A2(new_n432), .A3(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n494), .B(new_n500), .C1(new_n689), .C2(new_n690), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n632), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n619), .A3(new_n615), .A4(new_n614), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n432), .A2(new_n567), .A3(new_n615), .A4(new_n614), .ZN(new_n813));
  OAI22_X1  g627(.A1(new_n809), .A2(new_n812), .B1(new_n813), .B2(new_n674), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n792), .A3(new_n239), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n566), .B1(new_n632), .B2(new_n810), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n616), .A2(new_n641), .A3(new_n817), .A4(new_n640), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n617), .A2(KEYINPUT109), .A3(new_n676), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n806), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n666), .A2(new_n635), .A3(new_n670), .A4(new_n733), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n559), .A2(new_n658), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n695), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n746), .A2(new_n686), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n755), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n750), .B2(new_n751), .ZN(new_n826));
  AND4_X1   g640(.A1(KEYINPUT53), .A2(new_n805), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n805), .A2(new_n820), .A3(new_n826), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n827), .B1(KEYINPUT110), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n797), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n805), .A2(new_n820), .A3(new_n826), .A4(KEYINPUT53), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n797), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n796), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n830), .A2(KEYINPUT110), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n833), .A3(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n431), .A2(new_n721), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT112), .Z(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n365), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n789), .A2(new_n790), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n562), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n848), .A2(new_n735), .A3(new_n773), .A4(new_n777), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n781), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n773), .A2(new_n848), .A3(new_n777), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n735), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n722), .A2(new_n615), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n702), .A2(new_n703), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n704), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n849), .A2(new_n857), .A3(KEYINPUT50), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n745), .A2(new_n722), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT113), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n239), .A2(new_n562), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n631), .A2(new_n501), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n712), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n741), .A3(new_n852), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n843), .B1(new_n850), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n847), .A2(new_n781), .A3(new_n849), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(KEYINPUT51), .A3(new_n859), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(G952), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n871), .B(G953), .C1(new_n849), .C2(new_n729), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n712), .A2(new_n861), .A3(new_n862), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n634), .A2(new_n636), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n861), .A2(new_n362), .A3(new_n852), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT48), .B1(new_n877), .B2(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n870), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n838), .A2(new_n842), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n871), .A2(new_n218), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n771), .A2(new_n239), .A3(new_n365), .A4(new_n652), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT108), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n844), .B(KEYINPUT49), .Z(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n712), .A3(new_n857), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n218), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n830), .A2(new_n835), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n612), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n585), .A2(new_n587), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n592), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  XOR2_X1   g715(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n895), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n897), .A2(KEYINPUT116), .A3(new_n606), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT116), .B1(new_n897), .B2(new_n606), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n901), .ZN(G51));
  XOR2_X1   g723(.A(new_n763), .B(KEYINPUT57), .Z(new_n910));
  AOI21_X1  g724(.A(new_n797), .B1(new_n830), .B2(new_n835), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n837), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n428), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n897), .A2(new_n762), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT118), .B(new_n895), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n912), .B2(new_n428), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n894), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G54));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n897), .A2(new_n920), .A3(new_n498), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT119), .A3(new_n480), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n895), .C1(new_n480), .C2(new_n921), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT119), .B1(new_n921), .B2(new_n480), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G60));
  AOI22_X1  g739(.A1(new_n552), .A2(new_n623), .B1(new_n626), .B2(new_n551), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n926), .B(new_n929), .C1(new_n837), .C2(new_n911), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n895), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n834), .A2(new_n796), .A3(new_n837), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT111), .B1(new_n841), .B2(new_n836), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n926), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(G63));
  XNOR2_X1  g750(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n231), .A2(new_n224), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n896), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n223), .A2(new_n226), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n894), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n668), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G66));
  NOR3_X1   g760(.A1(new_n564), .A2(new_n590), .A3(new_n218), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n820), .B2(new_n218), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n899), .B1(G898), .B2(new_n218), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT122), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NAND3_X1  g765(.A1(new_n785), .A2(new_n752), .A3(new_n794), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n803), .A2(new_n717), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n362), .A2(new_n736), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n955), .B(new_n755), .C1(new_n768), .C2(new_n956), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n953), .B1(new_n952), .B2(new_n957), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n218), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n470), .A2(new_n471), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n335), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n955), .B(KEYINPUT62), .C1(new_n712), .C2(new_n707), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n713), .B2(new_n954), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n965), .A2(new_n967), .B1(new_n791), .B2(new_n793), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n745), .B(new_n699), .C1(new_n632), .C2(new_n810), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n362), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n785), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n785), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n968), .B(KEYINPUT125), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(G953), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n962), .B(KEYINPUT123), .Z(new_n979));
  OAI21_X1  g793(.A(new_n964), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n964), .B(new_n983), .C1(new_n978), .C2(new_n979), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n351), .B2(new_n708), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n840), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n958), .A2(new_n820), .A3(new_n959), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n987), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n336), .A2(new_n247), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n895), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n976), .A2(new_n820), .A3(new_n977), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n247), .B(new_n336), .C1(new_n995), .C2(new_n987), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n996), .ZN(G57));
endmodule


