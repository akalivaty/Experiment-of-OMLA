//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203));
  INV_X1    g002(.A(G57gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G64gat), .ZN(new_n205));
  INV_X1    g004(.A(G64gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G57gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT98), .ZN(new_n213));
  NOR2_X1   g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(KEYINPUT98), .B2(new_n212), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G71gat), .B(G78gat), .ZN(new_n217));
  AND4_X1   g016(.A1(KEYINPUT99), .A2(new_n208), .A3(new_n217), .A4(new_n210), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n209), .B1(new_n205), .B2(new_n207), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT99), .B1(new_n219), .B2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT101), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n208), .A2(new_n217), .A3(new_n210), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT99), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(KEYINPUT99), .A3(new_n217), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT101), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n216), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n203), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT16), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT94), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n233), .B(new_n235), .C1(new_n232), .C2(new_n231), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(KEYINPUT94), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n230), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT102), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(new_n242), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n202), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  INV_X1    g046(.A(new_n202), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n251));
  XNOR2_X1  g050(.A(G183gat), .B(G211gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  OR2_X1    g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n221), .A2(new_n203), .ZN(new_n255));
  NAND2_X1  g054(.A1(G231gat), .A2(G233gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT100), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n255), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n253), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n254), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G134gat), .B(G162gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(G29gat), .A2(G36gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(KEYINPUT14), .ZN(new_n269));
  INV_X1    g068(.A(new_n268), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT92), .B(G29gat), .ZN(new_n271));
  INV_X1    g070(.A(G36gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n273), .B2(KEYINPUT14), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT93), .ZN(new_n275));
  XOR2_X1   g074(.A(G43gat), .B(G50gat), .Z(new_n276));
  INV_X1    g075(.A(KEYINPUT15), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n280));
  INV_X1    g079(.A(new_n269), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n277), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n274), .B(new_n282), .C1(KEYINPUT93), .C2(new_n278), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT17), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n288), .A3(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT104), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT104), .A2(G99gat), .A3(G106gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G85gat), .ZN(new_n299));
  INV_X1    g098(.A(G92gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n296), .A2(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G99gat), .B(G106gat), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n303), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n305), .A2(new_n295), .A3(new_n298), .A4(new_n301), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT105), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n289), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n285), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n311), .A2(KEYINPUT106), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT106), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n316), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n309), .B(new_n319), .C1(new_n313), .C2(new_n314), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n318), .B1(new_n317), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n267), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n266), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT27), .B(G183gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n318), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NOR2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT26), .ZN(new_n336));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT65), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n336), .A2(new_n338), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n333), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n334), .B1(new_n333), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n343), .B2(new_n344), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  INV_X1    g146(.A(G183gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n318), .ZN(new_n349));
  NAND3_X1  g148(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(new_n350), .C1(G183gat), .C2(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n335), .A2(KEYINPUT23), .B1(KEYINPUT66), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n346), .A2(new_n351), .A3(new_n338), .A4(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(KEYINPUT66), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n357));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n358), .A2(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n359), .ZN(new_n367));
  INV_X1    g166(.A(new_n364), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(KEYINPUT68), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n357), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n357), .A3(new_n369), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  OAI22_X1  g171(.A1(new_n342), .A2(new_n356), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G227gat), .ZN(new_n374));
  INV_X1    g173(.A(G233gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n333), .A2(new_n339), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT67), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n333), .A2(new_n334), .A3(new_n339), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n372), .A2(new_n370), .ZN(new_n381));
  INV_X1    g180(.A(new_n355), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n354), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n373), .A2(new_n376), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G15gat), .B(G43gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n385), .B(KEYINPUT32), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT34), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n373), .A2(new_n384), .ZN(new_n397));
  INV_X1    g196(.A(new_n376), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT34), .B(new_n376), .C1(new_n373), .C2(new_n384), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n392), .A3(new_n394), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT71), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n394), .B2(new_n392), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT90), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT76), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT72), .B(G197gat), .Z(new_n421));
  INV_X1    g220(.A(G204gat), .ZN(new_n422));
  INV_X1    g221(.A(G211gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(new_n265), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n421), .A2(new_n422), .B1(KEYINPUT22), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n422), .B2(new_n421), .ZN(new_n426));
  XOR2_X1   g225(.A(G211gat), .B(G218gat), .Z(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n383), .A2(new_n377), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n356), .B1(new_n378), .B2(new_n379), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437));
  INV_X1    g236(.A(new_n431), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n380), .A2(new_n383), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT74), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n429), .B(new_n435), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n438), .B1(new_n436), .B2(KEYINPUT29), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n432), .A2(new_n431), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n429), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n440), .A2(KEYINPUT74), .A3(new_n431), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n434), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n429), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n420), .B(new_n444), .C1(new_n451), .C2(new_n443), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n431), .B1(new_n440), .B2(new_n433), .ZN(new_n457));
  INV_X1    g256(.A(new_n446), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n428), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n443), .B1(new_n442), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT75), .B1(new_n450), .B2(new_n429), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n419), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n452), .B2(new_n454), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n456), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G57gat), .B(G85gat), .Z(new_n466));
  XNOR2_X1  g265(.A(G1gat), .B(G29gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n471));
  XOR2_X1   g270(.A(G141gat), .B(G148gat), .Z(new_n472));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT2), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G155gat), .ZN(new_n476));
  INV_X1    g275(.A(G162gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n473), .ZN(new_n479));
  NOR2_X1   g278(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n475), .B(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT83), .B(new_n471), .C1(new_n381), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n365), .A2(new_n369), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT70), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n486), .B2(new_n371), .ZN(new_n487));
  INV_X1    g286(.A(new_n471), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n479), .A2(new_n480), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n475), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n485), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n483), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT81), .Z(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n482), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n485), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(KEYINPUT80), .A3(new_n499), .A4(new_n500), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n494), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n365), .A3(new_n369), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n496), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g312(.A(new_n496), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n492), .B2(new_n510), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n509), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n515), .B2(KEYINPUT85), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(KEYINPUT86), .C1(KEYINPUT85), .C2(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n506), .B1(new_n494), .B2(new_n505), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n508), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n488), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n503), .A2(new_n504), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT88), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n470), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n528), .B(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n494), .A2(new_n505), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n536), .A2(new_n507), .A3(new_n517), .A4(new_n520), .ZN(new_n537));
  INV_X1    g336(.A(new_n470), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n533), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT6), .B(new_n470), .C1(new_n523), .C2(new_n532), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n429), .A2(new_n433), .A3(new_n482), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n498), .A2(new_n433), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n428), .ZN(new_n546));
  AND2_X1   g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n500), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n482), .A2(new_n497), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n547), .ZN(new_n551));
  XOR2_X1   g350(.A(G78gat), .B(G106gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G22gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT31), .B(G50gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n551), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n415), .A2(new_n465), .A3(new_n543), .A4(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n541), .A2(new_n542), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n460), .A2(new_n419), .A3(new_n461), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT77), .B1(new_n561), .B2(KEYINPUT30), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT30), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n455), .A3(new_n462), .A4(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n403), .A2(new_n404), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n566), .A2(new_n559), .A3(new_n556), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n558), .A2(new_n559), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n411), .A2(new_n413), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n569), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n463), .A2(new_n464), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n543), .A2(new_n455), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n574), .B2(new_n556), .ZN(new_n575));
  OR3_X1    g374(.A1(new_n526), .A2(KEYINPUT39), .A3(new_n514), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n492), .A2(new_n510), .A3(new_n514), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT39), .B(new_n577), .C1(new_n526), .C2(new_n514), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n538), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT40), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n581), .A2(new_n533), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n585), .B(new_n444), .C1(new_n451), .C2(new_n443), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n435), .B1(new_n439), .B2(new_n441), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n588), .A3(new_n428), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT89), .B1(new_n450), .B2(new_n429), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n445), .A2(new_n429), .A3(new_n446), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n586), .B(new_n419), .C1(new_n592), .C2(new_n585), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n444), .B1(new_n451), .B2(new_n443), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(KEYINPUT37), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n460), .A2(new_n461), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n420), .B1(new_n597), .B2(new_n585), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n593), .A2(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n541), .A2(new_n542), .A3(new_n452), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n584), .B(new_n557), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n601), .ZN(new_n602));
  AOI211_X1 g401(.A(new_n263), .B(new_n329), .C1(new_n568), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  INV_X1    g403(.A(G197gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT11), .B(G169gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT97), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT18), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n240), .B1(new_n289), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n238), .A2(new_n614), .A3(new_n239), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n616), .A2(new_n288), .B1(new_n284), .B2(new_n285), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT96), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n613), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(new_n613), .C1(new_n615), .C2(new_n617), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n286), .A2(new_n240), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n286), .A2(new_n240), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n620), .B(KEYINPUT13), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n610), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n615), .A2(new_n617), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n612), .B1(new_n630), .B2(new_n620), .ZN(new_n631));
  INV_X1    g430(.A(new_n610), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n631), .A2(new_n632), .A3(new_n627), .A4(new_n623), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n307), .A2(new_n221), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n227), .A2(new_n304), .A3(new_n216), .A4(new_n306), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n306), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n222), .B2(new_n229), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(KEYINPUT107), .B(new_n641), .C1(new_n222), .C2(new_n229), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n636), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n637), .A2(new_n638), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n636), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n603), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n543), .B(KEYINPUT108), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT109), .B(G1gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1324gat));
  INV_X1    g459(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n564), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT16), .B(G8gat), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT110), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT110), .B(new_n667), .C1(new_n662), .C2(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(G8gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(G1325gat));
  AND3_X1   g469(.A1(new_n661), .A2(G15gat), .A3(new_n572), .ZN(new_n671));
  AOI21_X1  g470(.A(G15gat), .B1(new_n661), .B2(new_n415), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n656), .A2(new_n557), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n654), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n263), .A2(new_n634), .A3(new_n677), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n328), .B(new_n678), .C1(new_n568), .C2(new_n602), .ZN(new_n679));
  INV_X1    g478(.A(new_n657), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n271), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT111), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n575), .A2(new_n601), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT90), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n557), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n559), .B1(new_n691), .B2(new_n574), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n565), .A2(new_n567), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n329), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n328), .B1(new_n568), .B2(new_n602), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n678), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n680), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n684), .B(new_n687), .C1(new_n271), .C2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n678), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n568), .A2(new_n602), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n698), .B1(new_n705), .B2(new_n329), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT44), .B(new_n328), .C1(new_n568), .C2(new_n602), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n708), .B2(new_n465), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n697), .A2(new_n272), .A3(new_n564), .A4(new_n704), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT112), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1329gat));
  OAI211_X1 g516(.A(new_n572), .B(new_n704), .C1(new_n706), .C2(new_n707), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n679), .A2(new_n720), .A3(new_n415), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1330gat));
  NAND2_X1  g523(.A1(new_n556), .A2(G50gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n695), .A2(new_n557), .A3(new_n678), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n708), .A2(new_n725), .B1(G50gat), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n677), .A2(new_n634), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n603), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n657), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n204), .ZN(G1332gat));
  AOI21_X1  g531(.A(new_n465), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n603), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT113), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  INV_X1    g536(.A(new_n415), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n730), .A2(G71gat), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n740));
  INV_X1    g539(.A(new_n572), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n740), .B1(new_n739), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n557), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g546(.A1(new_n262), .A2(new_n634), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n654), .B(new_n748), .C1(new_n706), .C2(new_n707), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n657), .ZN(new_n750));
  AND4_X1   g549(.A1(KEYINPUT51), .A2(new_n705), .A3(new_n329), .A4(new_n748), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT51), .B1(new_n697), .B2(new_n748), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n680), .A2(new_n299), .A3(new_n654), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT114), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(G1336gat));
  OAI211_X1 g555(.A(new_n564), .B(new_n654), .C1(new_n751), .C2(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n300), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n748), .A2(new_n654), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n696), .B2(new_n699), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n465), .A2(new_n300), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n758), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n758), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1337gat));
  OR4_X1    g567(.A1(G99gat), .A2(new_n753), .A3(new_n738), .A4(new_n677), .ZN(new_n769));
  OAI21_X1  g568(.A(G99gat), .B1(new_n749), .B2(new_n741), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  OAI21_X1  g570(.A(G106gat), .B1(new_n749), .B2(new_n557), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n557), .A2(G106gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n654), .B(new_n773), .C1(new_n751), .C2(new_n752), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n774), .B2(KEYINPUT116), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n772), .B(new_n774), .C1(KEYINPUT116), .C2(new_n776), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1339gat));
  OR3_X1    g579(.A1(new_n644), .A2(new_n636), .A3(new_n645), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n783), .B(new_n636), .C1(new_n644), .C2(new_n645), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n784), .A2(KEYINPUT117), .A3(new_n651), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT117), .B1(new_n784), .B2(new_n651), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT55), .B(new_n782), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n789), .A2(new_n634), .A3(new_n652), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n618), .A2(new_n621), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n626), .B1(new_n624), .B2(new_n625), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n608), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n654), .A2(new_n633), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n791), .A2(KEYINPUT118), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT118), .B1(new_n791), .B2(new_n795), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(new_n329), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n789), .A2(new_n652), .A3(new_n790), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n633), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n328), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n263), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n634), .A2(new_n654), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n262), .A2(new_n328), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n691), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n657), .A2(new_n564), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n635), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n556), .B(new_n566), .C1(new_n802), .C2(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n635), .A2(G113gat), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT119), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n808), .B1(new_n810), .B2(new_n812), .ZN(G1340gat));
  OAI21_X1  g612(.A(G120gat), .B1(new_n807), .B2(new_n677), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n677), .A2(G120gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n810), .B2(new_n815), .ZN(G1341gat));
  INV_X1    g615(.A(new_n810), .ZN(new_n817));
  AOI21_X1  g616(.A(G127gat), .B1(new_n817), .B2(new_n262), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n805), .A2(G127gat), .A3(new_n262), .A4(new_n806), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(KEYINPUT120), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(KEYINPUT120), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(G1342gat));
  NOR4_X1   g621(.A1(new_n657), .A2(G134gat), .A3(new_n564), .A4(new_n328), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n809), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT56), .Z(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n807), .B2(new_n328), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1343gat));
  NOR2_X1   g626(.A1(new_n657), .A2(new_n572), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n465), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n329), .B1(new_n791), .B2(new_n795), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n263), .B1(new_n830), .B2(new_n801), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n557), .B1(new_n831), .B2(new_n804), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT57), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT121), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n557), .B1(new_n802), .B2(new_n804), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n829), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n634), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G141gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  INV_X1    g641(.A(new_n829), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n835), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(G141gat), .A3(new_n635), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(G141gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n839), .B2(new_n634), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT58), .B1(new_n849), .B2(new_n845), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(G1344gat));
  INV_X1    g650(.A(new_n844), .ZN(new_n852));
  INV_X1    g651(.A(G148gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n654), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT59), .B(new_n853), .C1(new_n839), .C2(new_n654), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n791), .A2(new_n795), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n329), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n791), .A2(KEYINPUT118), .A3(new_n795), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n801), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n804), .B1(new_n861), .B2(new_n262), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n556), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT122), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT57), .A4(new_n556), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT123), .B1(new_n832), .B2(KEYINPUT57), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n799), .A2(new_n328), .A3(new_n800), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n857), .A2(new_n328), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n262), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n804), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n556), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n837), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n654), .A3(new_n843), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n856), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n854), .B1(new_n855), .B2(new_n877), .ZN(G1345gat));
  AOI21_X1  g677(.A(G155gat), .B1(new_n852), .B2(new_n262), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n263), .A2(new_n476), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n839), .B2(new_n880), .ZN(G1346gat));
  NAND2_X1  g680(.A1(new_n839), .A2(new_n329), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G162gat), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n828), .A2(new_n477), .A3(new_n465), .A4(new_n329), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n836), .B2(new_n884), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n680), .A2(new_n465), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n809), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(G169gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n634), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n805), .A2(new_n886), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n805), .A2(new_n886), .A3(KEYINPUT124), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n634), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n890), .B1(new_n896), .B2(new_n889), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n888), .B2(new_n654), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n654), .A2(G176gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n262), .A3(new_n894), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G183gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n888), .A2(new_n330), .A3(new_n262), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n318), .A3(new_n329), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n895), .A2(new_n329), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(G190gat), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT61), .B(new_n318), .C1(new_n895), .C2(new_n329), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  NOR3_X1   g710(.A1(new_n680), .A2(new_n465), .A3(new_n572), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n835), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(G197gat), .A3(new_n635), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n875), .A2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n634), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(new_n605), .ZN(G1352gat));
  INV_X1    g718(.A(new_n913), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n422), .A3(new_n654), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n921), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n875), .A2(new_n654), .A3(new_n912), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G204gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(new_n921), .B2(KEYINPUT62), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n922), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n920), .A2(new_n423), .A3(new_n262), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n865), .B1(new_n835), .B2(KEYINPUT57), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n262), .B(new_n912), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n875), .A2(new_n933), .A3(new_n262), .A4(new_n912), .ZN(new_n934));
  AND4_X1   g733(.A1(KEYINPUT63), .A2(new_n932), .A3(G211gat), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n423), .B1(new_n931), .B2(KEYINPUT127), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n936), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n928), .B1(new_n935), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n920), .B2(new_n329), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n328), .A2(new_n265), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n916), .B2(new_n940), .ZN(G1355gat));
endmodule


