//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n591, new_n593, new_n594, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n464), .B2(new_n465), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n480), .B1(new_n468), .B2(G136), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n469), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .A4(new_n469), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n487), .A2(new_n489), .A3(new_n490), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  OR2_X1    g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(G88), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n502), .A2(new_n508), .ZN(G166));
  INV_X1    g084(.A(new_n506), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT7), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(KEYINPUT7), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G51), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n497), .A2(new_n498), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n503), .A2(G89), .ZN(new_n517));
  NAND2_X1  g092(.A1(G63), .A2(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G168));
  AOI22_X1  g095(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT71), .B(G90), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n504), .A2(new_n523), .B1(new_n506), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G171));
  AOI22_X1  g101(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n501), .ZN(new_n528));
  INV_X1    g103(.A(G81), .ZN(new_n529));
  INV_X1    g104(.A(G43), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n504), .A2(new_n529), .B1(new_n506), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G860), .ZN(G153));
  AND3_X1   g108(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G36), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n534), .A2(new_n538), .ZN(G188));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n503), .A2(new_n540), .A3(G53), .A4(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT9), .ZN(new_n542));
  NAND2_X1  g117(.A1(G78), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n516), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n504), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G651), .B1(new_n546), .B2(G91), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(G299));
  INV_X1    g123(.A(G171), .ZN(G301));
  INV_X1    g124(.A(G168), .ZN(G286));
  INV_X1    g125(.A(G166), .ZN(G303));
  OAI21_X1  g126(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n499), .A2(new_n503), .A3(G87), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n503), .A2(G49), .A3(G543), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(G288));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n497), .B2(new_n498), .ZN(new_n563));
  AND2_X1   g138(.A1(G73), .A2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n546), .B2(G86), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n503), .A2(KEYINPUT75), .A3(G48), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n566), .A2(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(G85), .A2(new_n546), .B1(new_n510), .B2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n501), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n499), .A2(new_n503), .A3(G92), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n516), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n510), .B2(G54), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n577), .B1(new_n584), .B2(G868), .ZN(G284));
  OAI21_X1  g160(.A(new_n577), .B1(new_n584), .B2(G868), .ZN(G321));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(G299), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n587), .B2(G168), .ZN(G297));
  OAI21_X1  g164(.A(new_n588), .B1(new_n587), .B2(G168), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n591), .B2(G860), .ZN(G148));
  NAND2_X1  g167(.A1(new_n584), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n532), .ZN(G323));
  XNOR2_X1  g170(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g171(.A1(new_n468), .A2(G2104), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT12), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT13), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(G2100), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n480), .A2(G123), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT77), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n468), .A2(G135), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT76), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n469), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n602), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G2096), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(G2096), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n600), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g186(.A(G2427), .B(G2438), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2430), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT15), .B(G2435), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(KEYINPUT14), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G1341), .B(G1348), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2443), .B(G2446), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(G2451), .B(G2454), .Z(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(G14), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(G401));
  XNOR2_X1  g203(.A(G2072), .B(G2078), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT17), .ZN(new_n630));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2067), .B(G2678), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT81), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n631), .A2(new_n629), .A3(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n630), .A2(new_n633), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(new_n632), .C1(new_n629), .C2(new_n633), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2096), .B(G2100), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(G227));
  XNOR2_X1  g218(.A(G1956), .B(G2474), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1961), .B(G1966), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT82), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  OR3_X1    g227(.A1(new_n644), .A2(new_n652), .A3(KEYINPUT82), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT20), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n644), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  MUX2_X1   g232(.A(new_n657), .B(new_n656), .S(new_n651), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(new_n662), .B2(new_n666), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n662), .A2(new_n666), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n667), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n676), .B2(new_n669), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G29), .A2(G35), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(G162), .B2(G29), .ZN(new_n680));
  INV_X1    g255(.A(G2090), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT25), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n468), .A2(G139), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT91), .Z(new_n690));
  AND2_X1   g265(.A1(new_n488), .A2(G127), .ZN(new_n691));
  AND2_X1   g266(.A1(G115), .A2(G2104), .ZN(new_n692));
  OAI21_X1  g267(.A(G2105), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G33), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2072), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT30), .B(G28), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  OR2_X1    g273(.A1(KEYINPUT31), .A2(G11), .ZN(new_n699));
  NAND2_X1  g274(.A1(KEYINPUT31), .A2(G11), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n607), .B2(new_n698), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  NOR3_X1   g278(.A1(new_n684), .A2(new_n696), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n468), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n480), .A2(G129), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n470), .A2(G105), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n698), .ZN(new_n713));
  MUX2_X1   g288(.A(new_n706), .B(KEYINPUT92), .S(new_n713), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G5), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G171), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n724), .B2(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(KEYINPUT24), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n472), .B2(new_n698), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n721), .A2(new_n722), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n717), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT94), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n532), .B2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT89), .B(G1341), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n734), .B1(new_n722), .B2(new_n721), .C1(new_n723), .C2(new_n727), .ZN(new_n735));
  NOR2_X1   g310(.A1(G4), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n584), .B2(G16), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT88), .B(G1348), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n698), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n468), .A2(G140), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT90), .Z(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n744));
  INV_X1    g319(.A(G116), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G2105), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n480), .B2(G128), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n718), .A2(G20), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT23), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G299), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n735), .A2(new_n739), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n718), .ZN(new_n759));
  INV_X1    g334(.A(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n698), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n761), .B(new_n765), .C1(new_n716), .C2(new_n714), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n682), .B2(new_n683), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n704), .A2(new_n730), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n468), .A2(G131), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT84), .Z(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G107), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT85), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n480), .A2(G119), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n770), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G25), .B(new_n776), .S(G29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT86), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XOR2_X1   g356(.A(KEYINPUT32), .B(G1981), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n718), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n718), .A2(G23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n555), .B2(new_n718), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n783), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  MUX2_X1   g368(.A(G24), .B(G290), .S(G16), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT87), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1986), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n780), .A2(new_n793), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT36), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT36), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n768), .B1(new_n799), .B2(new_n800), .ZN(G311));
  XNOR2_X1  g376(.A(G311), .B(KEYINPUT96), .ZN(G150));
  NAND2_X1  g377(.A1(new_n584), .A2(G559), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n501), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n504), .A2(new_n808), .B1(new_n506), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n532), .A2(new_n811), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n528), .A2(new_n531), .B1(new_n807), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n805), .B(new_n814), .Z(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(G860), .ZN(new_n818));
  INV_X1    g393(.A(new_n811), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  OR2_X1    g397(.A1(new_n818), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n607), .B(new_n472), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n487), .A2(new_n489), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n490), .A2(new_n494), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n490), .A2(KEYINPUT99), .A3(new_n494), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n748), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n694), .A2(new_n712), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n480), .A2(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n468), .A2(G142), .ZN(new_n836));
  OR2_X1    g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n712), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n690), .A2(new_n693), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n834), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n833), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n834), .A2(new_n841), .ZN(new_n845));
  INV_X1    g420(.A(new_n839), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n832), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n776), .B(new_n598), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT100), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n844), .B2(new_n849), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n825), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n844), .A2(new_n849), .ZN(new_n855));
  INV_X1    g430(.A(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n851), .A4(new_n824), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G162), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  INV_X1    g436(.A(G162), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n854), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(G395));
  XNOR2_X1  g441(.A(new_n584), .B(G299), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT41), .Z(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n593), .B(new_n814), .Z(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n873), .A2(KEYINPUT42), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n555), .B(KEYINPUT103), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(G290), .B(G166), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n873), .B2(new_n874), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n875), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n875), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n811), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n811), .ZN(G331));
  NAND2_X1  g461(.A1(G171), .A2(KEYINPUT105), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n814), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  AOI21_X1  g464(.A(G168), .B1(G301), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n868), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n867), .A3(new_n892), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n880), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n861), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n880), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n861), .A4(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(KEYINPUT106), .A3(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n903), .ZN(G397));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n490), .A2(KEYINPUT99), .A3(new_n494), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT99), .B1(new_n490), .B2(new_n494), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n914), .B2(new_n826), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(G1996), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT108), .B1(new_n919), .B2(new_n840), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n748), .B(new_n750), .ZN(new_n921));
  INV_X1    g496(.A(G1996), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n840), .ZN(new_n923));
  INV_X1    g498(.A(new_n918), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(KEYINPUT108), .A3(new_n840), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n776), .B(new_n779), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n918), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n918), .A2(G1986), .A3(G290), .ZN(new_n930));
  AND2_X1   g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT107), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT109), .ZN(new_n935));
  INV_X1    g510(.A(G8), .ZN(new_n936));
  NOR2_X1   g511(.A1(G166), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n487), .A2(new_n489), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n913), .B2(new_n912), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(new_n911), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n829), .A2(new_n830), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n946), .B2(new_n941), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT113), .B(new_n917), .C1(new_n947), .C2(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n495), .A2(new_n911), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n945), .A2(new_n681), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n944), .B1(new_n949), .B2(new_n916), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT45), .B(new_n911), .C1(new_n914), .C2(new_n826), .ZN(new_n954));
  AOI21_X1  g529(.A(G1971), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n938), .B1(new_n957), .B2(G8), .ZN(new_n958));
  INV_X1    g533(.A(G1981), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n546), .A2(G86), .ZN(new_n960));
  OAI21_X1  g535(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n571), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n566), .A2(new_n964), .A3(new_n959), .A4(new_n571), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G305), .A2(G1981), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(KEYINPUT49), .A3(new_n967), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n942), .A2(new_n911), .A3(new_n917), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n555), .A2(G1976), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(G8), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(KEYINPUT52), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n560), .B2(G1976), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n944), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n940), .B(new_n911), .C1(new_n914), .C2(new_n826), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G2090), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n938), .B(G8), .C1(new_n986), .C2(new_n955), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n975), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n958), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n917), .B1(new_n947), .B2(KEYINPUT45), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n495), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n911), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G2078), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OR3_X1    g573(.A1(new_n990), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n953), .A2(new_n954), .A3(new_n764), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n1000), .A2(new_n996), .B1(new_n985), .B2(new_n722), .ZN(new_n1001));
  AOI21_X1  g576(.A(G301), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n760), .B1(new_n990), .B2(new_n995), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n983), .A2(new_n984), .A3(new_n723), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(G168), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(G168), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1003), .B1(KEYINPUT62), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(KEYINPUT62), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G286), .A2(new_n936), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n989), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n1019));
  INV_X1    g594(.A(new_n975), .ZN(new_n1020));
  OR2_X1    g595(.A1(G288), .A2(G1976), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1019), .B(new_n966), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n973), .B1(new_n968), .B2(new_n969), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(new_n971), .ZN(new_n1024));
  INV_X1    g599(.A(new_n966), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT112), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n973), .B(KEYINPUT111), .Z(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n986), .A2(new_n955), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n936), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(new_n938), .A3(new_n975), .A4(new_n982), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1016), .B(new_n1017), .C1(new_n1030), .C2(new_n938), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT63), .B1(new_n1032), .B2(new_n988), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1018), .A2(new_n1028), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n948), .A2(new_n951), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT50), .B1(new_n831), .B2(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n917), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n755), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n542), .B2(KEYINPUT115), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G299), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n542), .B(new_n547), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n953), .A2(new_n954), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1348), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n985), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n915), .A2(new_n944), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n750), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1051), .A3(KEYINPUT116), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1348), .B1(new_n983), .B2(new_n984), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n915), .A2(G2067), .A3(new_n944), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1047), .A2(new_n584), .A3(new_n1052), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n944), .B1(new_n915), .B2(KEYINPUT50), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n950), .B1(new_n1058), .B2(KEYINPUT113), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1956), .B1(new_n1059), .B2(new_n945), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1046), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1042), .A2(KEYINPUT117), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1042), .A2(KEYINPUT117), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1060), .A2(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1052), .A2(new_n1066), .A3(new_n1056), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n584), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1069), .B2(new_n584), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n584), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT119), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1070), .A3(new_n584), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1067), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1047), .A2(KEYINPUT118), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1038), .A2(new_n1080), .A3(new_n1042), .A4(new_n1046), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(KEYINPUT61), .A3(new_n1081), .A4(new_n1064), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1047), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1042), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1043), .A2(G1996), .B1(new_n1050), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n532), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT59), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1065), .B1(new_n1078), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n985), .B2(new_n722), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT120), .B(G1961), .C1(new_n983), .C2(new_n984), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1000), .A2(new_n996), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n915), .A2(new_n916), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(new_n917), .A3(new_n954), .A4(new_n997), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1097), .A2(G171), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1093), .B1(new_n1102), .B2(new_n1002), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1012), .A2(new_n989), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n999), .A2(G301), .A3(new_n1001), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT121), .ZN(new_n1106));
  OAI21_X1  g681(.A(G171), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n999), .A2(new_n1001), .A3(new_n1108), .A4(G301), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT54), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT122), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1107), .A2(KEYINPUT54), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1109), .A4(new_n1106), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1104), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1034), .B1(new_n1092), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1014), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g693(.A(KEYINPUT123), .B(new_n1034), .C1(new_n1092), .C2(new_n1115), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n935), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n779), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n776), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n927), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n743), .A2(new_n750), .A3(new_n747), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n918), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n918), .B1(new_n921), .B2(new_n840), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT46), .B1(new_n918), .B2(G1996), .ZN(new_n1130));
  OR3_X1    g705(.A1(new_n918), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n930), .B(KEYINPUT48), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n929), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1127), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1120), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g713(.A1(G227), .A2(new_n458), .ZN(new_n1140));
  OAI211_X1 g714(.A(new_n627), .B(new_n1140), .C1(new_n674), .C2(new_n677), .ZN(new_n1141));
  AOI21_X1  g715(.A(new_n1141), .B1(new_n899), .B2(new_n902), .ZN(new_n1142));
  AND3_X1   g716(.A1(new_n1142), .A2(new_n864), .A3(KEYINPUT126), .ZN(new_n1143));
  AOI21_X1  g717(.A(KEYINPUT126), .B1(new_n1142), .B2(new_n864), .ZN(new_n1144));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n1144), .ZN(G308));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n864), .ZN(G225));
endmodule


