//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR3_X1   g042(.A1(new_n466), .A2(new_n467), .A3(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G101), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n469), .B1(new_n462), .B2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT66), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n480), .B(new_n483), .C1(G136), .C2(new_n464), .ZN(G162));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(new_n490), .B1(new_n481), .B2(G126), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n469), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n473), .A2(new_n496), .A3(G138), .A4(new_n469), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AND3_X1   g079(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT5), .B1(KEYINPUT68), .B2(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(G62), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n507), .B2(KEYINPUT69), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(G62), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(G50), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n505), .A2(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n501), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT68), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n503), .B1(new_n524), .B2(new_n509), .ZN(new_n525));
  INV_X1    g100(.A(new_n510), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n517), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(KEYINPUT70), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n518), .A2(new_n529), .ZN(G166));
  NAND2_X1  g105(.A1(new_n522), .A2(new_n523), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(G89), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(G51), .A3(G543), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n515), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(G64), .B1(new_n505), .B2(new_n506), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n502), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT71), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n522), .B2(new_n523), .ZN(new_n549));
  INV_X1    g124(.A(new_n545), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n532), .A2(G52), .A3(G543), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n531), .A2(G90), .A3(new_n532), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n547), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n502), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n515), .A2(new_n559), .B1(new_n541), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT72), .Z(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT73), .ZN(G188));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n541), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n532), .A2(new_n572), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n522), .B2(new_n523), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n515), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G91), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n574), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n584));
  NOR2_X1   g159(.A1(G166), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT74), .B1(new_n518), .B2(new_n529), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G303));
  NAND2_X1  g162(.A1(new_n579), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(new_n541), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G49), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(G288));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n522), .B2(new_n523), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n595));
  INV_X1    g170(.A(G73), .ZN(new_n596));
  INV_X1    g171(.A(G543), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(G61), .B1(new_n505), .B2(new_n506), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  INV_X1    g177(.A(G48), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n515), .A2(new_n602), .B1(new_n541), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  NAND3_X1  g181(.A1(new_n531), .A2(G85), .A3(new_n532), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT76), .B(G47), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n532), .A2(new_n608), .A3(G543), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n607), .B(new_n609), .C1(new_n610), .C2(new_n502), .ZN(G290));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n612));
  OAI21_X1  g187(.A(G66), .B1(new_n505), .B2(new_n506), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n502), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n532), .A2(G54), .A3(G543), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n531), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  OAI211_X1 g194(.A(KEYINPUT77), .B(new_n616), .C1(new_n619), .C2(new_n502), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n515), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(G301), .B(new_n625), .S(new_n626), .Z(G284));
  MUX2_X1   g202(.A(G301), .B(new_n625), .S(new_n626), .Z(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n581), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(new_n625), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(G860), .B2(new_n633), .ZN(G148));
  OAI21_X1  g209(.A(KEYINPUT80), .B1(new_n562), .B2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  MUX2_X1   g213(.A(KEYINPUT80), .B(new_n635), .S(new_n638), .Z(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g215(.A1(new_n468), .A2(new_n470), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n473), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n464), .A2(G135), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n481), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n469), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT82), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT14), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(KEYINPUT83), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(KEYINPUT83), .ZN(new_n662));
  OAI22_X1  g237(.A1(new_n661), .A2(new_n662), .B1(new_n656), .B2(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(KEYINPUT84), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(KEYINPUT84), .A3(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n681), .B2(new_n678), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(KEYINPUT20), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n697), .B1(new_n694), .B2(new_n698), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1981), .B(G1986), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n706), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n709), .B1(new_n707), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n691), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n690), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n720), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(G1971), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G23), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT90), .Z(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G288), .B2(new_n720), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n720), .A2(G6), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n596), .A2(new_n597), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n599), .B2(KEYINPUT75), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n594), .A2(new_n595), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n502), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n604), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(new_n720), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT32), .B(G1981), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT89), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n723), .A2(new_n724), .A3(new_n729), .A4(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n607), .A2(new_n609), .ZN(new_n743));
  OAI21_X1  g318(.A(G60), .B1(new_n505), .B2(new_n506), .ZN(new_n744));
  NAND2_X1  g319(.A1(G72), .A2(G543), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n502), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(new_n720), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n720), .B2(G24), .ZN(new_n749));
  INV_X1    g324(.A(G1986), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n464), .A2(G131), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n481), .A2(G119), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n469), .A2(G107), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G25), .B(new_n756), .S(G29), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT35), .B(G1991), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n757), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n749), .A2(new_n750), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n741), .A2(new_n742), .A3(new_n751), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT36), .Z(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(G164), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G27), .B2(new_n765), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n720), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n720), .B2(G21), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n768), .A2(G2078), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n765), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n765), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n772), .B1(new_n769), .B2(new_n771), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n774), .A2(new_n778), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT30), .B(G28), .ZN(new_n781));
  OR2_X1    g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n765), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n652), .B2(new_n765), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n765), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n464), .A2(G140), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n481), .A2(G128), .ZN(new_n790));
  OR2_X1    g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n788), .B1(new_n794), .B2(new_n765), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G2078), .B2(new_n768), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n779), .A2(new_n780), .A3(new_n786), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n720), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n632), .B2(new_n720), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n804), .A2(G5), .A3(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(G5), .B2(G16), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(G301), .C2(new_n720), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n720), .A2(G20), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT23), .Z(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G105), .B2(new_n641), .ZN(new_n819));
  AOI22_X1  g394(.A1(G129), .A2(new_n481), .B1(new_n464), .B2(G141), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n765), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n765), .B2(G32), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT27), .B(G1996), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(KEYINPUT24), .A2(G34), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n765), .B1(KEYINPUT24), .B2(G34), .ZN(new_n828));
  OAI22_X1  g403(.A1(G160), .A2(new_n765), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n826), .B1(G2084), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(G2084), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n824), .B2(new_n825), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n765), .A2(G33), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n464), .A2(G139), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT92), .Z(new_n835));
  NAND3_X1  g410(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT91), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT25), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n473), .A2(G127), .ZN(new_n839));
  INV_X1    g414(.A(G115), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n467), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G2105), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n835), .B(new_n838), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n833), .B1(new_n845), .B2(G29), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(G2072), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n720), .A2(G19), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n562), .B2(new_n720), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(G1341), .Z(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n847), .B2(G2072), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n830), .A2(new_n832), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n799), .A2(new_n803), .A3(new_n815), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n764), .A2(new_n854), .ZN(G311));
  INV_X1    g430(.A(G311), .ZN(G150));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n522), .B2(new_n523), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(G67), .B1(new_n505), .B2(new_n506), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n859), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(G651), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT99), .ZN(new_n866));
  INV_X1    g441(.A(G93), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n515), .A2(new_n867), .B1(new_n541), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT100), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n871), .B1(new_n541), .B2(new_n868), .C1(new_n515), .C2(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n861), .A2(new_n874), .A3(G651), .A4(new_n864), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n562), .A2(KEYINPUT101), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n558), .B2(new_n561), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(KEYINPUT99), .A2(new_n865), .B1(new_n870), .B2(new_n872), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(KEYINPUT101), .A3(new_n562), .A4(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT38), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n632), .A2(G559), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n884), .B(new_n885), .Z(new_n886));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g462(.A(G860), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n876), .A2(G860), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT37), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G145));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n821), .B1(new_n845), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n845), .A2(new_n893), .A3(new_n821), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n464), .A2(G142), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n481), .A2(G130), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n469), .A2(G118), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n897), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n756), .B(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n895), .B2(new_n896), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT102), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT102), .B1(new_n495), .B2(new_n497), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n491), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n794), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n644), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n904), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G160), .B(new_n652), .ZN(new_n914));
  XNOR2_X1  g489(.A(G162), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n915), .B2(new_n913), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g493(.A(new_n883), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n637), .B(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n621), .A2(new_n581), .A3(new_n624), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n581), .B1(new_n621), .B2(new_n624), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n921), .B2(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n625), .A2(G299), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n621), .A2(new_n581), .A3(new_n624), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n925), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n601), .A2(new_n605), .A3(G290), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n747), .B1(new_n734), .B2(new_n604), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n518), .A2(new_n529), .A3(G288), .ZN(new_n938));
  AOI21_X1  g513(.A(G288), .B1(new_n518), .B2(new_n529), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G288), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT70), .B1(new_n527), .B2(new_n528), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n510), .A3(new_n503), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n501), .B(new_n517), .C1(new_n944), .C2(G651), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n518), .A2(new_n529), .A3(G288), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n935), .A2(new_n936), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n940), .A2(KEYINPUT105), .A3(new_n949), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT105), .B1(new_n940), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  MUX2_X1   g529(.A(new_n950), .B(new_n954), .S(KEYINPUT42), .Z(new_n955));
  AND2_X1   g530(.A1(new_n934), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n934), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n876), .A2(new_n626), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n959), .ZN(G331));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n547), .A2(new_n555), .A3(G286), .ZN(new_n963));
  AOI21_X1  g538(.A(G286), .B1(new_n547), .B2(new_n555), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n880), .A2(new_n965), .A3(new_n882), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n880), .B2(new_n882), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n933), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n883), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n880), .A2(new_n965), .A3(new_n882), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n923), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(new_n972), .A3(KEYINPUT106), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n970), .A2(new_n923), .A3(new_n974), .A4(new_n971), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n953), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n962), .B1(new_n976), .B2(KEYINPUT107), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n978), .B(new_n953), .C1(new_n973), .C2(new_n975), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n953), .A3(new_n975), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT108), .B1(new_n923), .B2(new_n926), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n930), .B2(new_n923), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n984), .B(new_n985), .C1(new_n966), .C2(new_n967), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n954), .B1(new_n986), .B2(new_n972), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NOR4_X1   g563(.A1(new_n977), .A2(new_n979), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT44), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n980), .B2(new_n981), .ZN(new_n992));
  NOR4_X1   g567(.A1(new_n977), .A2(new_n979), .A3(new_n987), .A4(KEYINPUT43), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT126), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT45), .B1(new_n908), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(G40), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n472), .A2(new_n476), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OR3_X1    g576(.A1(new_n1001), .A2(KEYINPUT112), .A3(G1996), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT112), .B1(new_n1001), .B2(G1996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n996), .B1(new_n1004), .B2(KEYINPUT46), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(KEYINPUT126), .A3(new_n1006), .A4(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n793), .B(G2067), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT113), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n1011), .B2(new_n822), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n1004), .B2(KEYINPUT46), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1008), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n821), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n821), .A2(G1996), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n756), .A2(new_n759), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(new_n796), .B2(new_n794), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n756), .B(new_n758), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1001), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1001), .A2(G1986), .A3(G290), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1022), .A2(new_n1001), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT127), .B1(new_n1016), .B2(new_n1029), .ZN(new_n1030));
  NOR4_X1   g605(.A1(new_n1028), .A2(new_n1017), .A3(new_n1019), .A4(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n794), .A2(new_n796), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1001), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT127), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1036), .B(new_n1037), .C1(new_n1015), .C2(new_n1014), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n908), .A2(new_n997), .A3(new_n1000), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  OR2_X1    g616(.A1(G305), .A2(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G305), .A2(G1981), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n941), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1042), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1041), .B1(new_n1051), .B2(KEYINPUT117), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1053), .A3(new_n1042), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT115), .B(KEYINPUT116), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G303), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  NAND3_X1  g638(.A1(G303), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n474), .A2(new_n475), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G2105), .ZN(new_n1066));
  INV_X1    g641(.A(new_n999), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n471), .A3(new_n465), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n499), .A2(new_n997), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT45), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n908), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1971), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1068), .B1(new_n1069), .B2(KEYINPUT50), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n908), .A2(new_n997), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(G2090), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1062), .A2(G8), .A3(new_n1064), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1040), .B(G8), .C1(new_n1049), .C2(G288), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n941), .A2(G1976), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1083), .A2(KEYINPUT52), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(KEYINPUT52), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1048), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1052), .A2(new_n1054), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1077), .B1(new_n908), .B2(new_n997), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1000), .B1(new_n1069), .B2(KEYINPUT50), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1075), .B1(new_n1091), .B2(G2090), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1064), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1063), .B1(G303), .B2(new_n1059), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1000), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n769), .B1(new_n998), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(G2084), .B2(new_n1079), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1099), .A2(G8), .A3(G168), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(new_n1081), .A3(new_n1087), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1100), .A2(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1080), .A2(G8), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1106));
  AND4_X1   g681(.A1(new_n1081), .A2(new_n1104), .A3(new_n1087), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1088), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1099), .B2(G286), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1079), .A2(G2084), .ZN(new_n1110));
  AOI21_X1  g685(.A(G168), .B1(new_n1110), .B2(new_n1098), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(G8), .C1(new_n1099), .C2(G286), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n998), .A2(new_n1097), .ZN(new_n1117));
  INV_X1    g692(.A(G2078), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1121), .A3(new_n1118), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(KEYINPUT53), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1073), .B2(G2078), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1079), .A2(new_n808), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G301), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1112), .A2(new_n1129), .A3(new_n1114), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1116), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n581), .B(KEYINPUT57), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n813), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1071), .A2(new_n1072), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1040), .A2(G2067), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n802), .B2(new_n1079), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(new_n625), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1133), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1137), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1133), .A2(KEYINPUT118), .A3(new_n1135), .A4(new_n1132), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(KEYINPUT61), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1040), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1073), .B2(G1996), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n562), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1154), .A3(new_n562), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1148), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1138), .B(KEYINPUT60), .C1(new_n1160), .C2(G1348), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(KEYINPUT119), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1161), .A2(KEYINPUT119), .A3(new_n625), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n625), .B1(new_n1161), .B2(KEYINPUT119), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1140), .A2(KEYINPUT60), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1144), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1065), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n474), .A2(KEYINPUT121), .A3(new_n475), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(G2105), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(G40), .A3(new_n471), .A4(new_n465), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AND2_X1   g751(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1177));
  NOR2_X1   g752(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT53), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1180));
  INV_X1    g755(.A(new_n998), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1176), .A2(new_n1180), .A3(new_n1181), .A4(new_n1072), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(G171), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1169), .B1(new_n1128), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(G171), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT125), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1123), .A2(G301), .A3(new_n1127), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1183), .A2(new_n1189), .A3(G171), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT54), .A4(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1185), .A2(new_n1191), .A3(new_n1115), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1131), .B1(new_n1168), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1096), .A2(new_n1081), .A3(new_n1087), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT124), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1108), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT110), .B1(new_n747), .B2(new_n750), .ZN(new_n1197));
  NAND2_X1  g772(.A1(G290), .A2(G1986), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1001), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT111), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1020), .A2(new_n1025), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1039), .B1(new_n1196), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g778(.A1(new_n992), .A2(new_n993), .ZN(new_n1205));
  OR2_X1    g779(.A1(new_n671), .A2(new_n672), .ZN(new_n1206));
  AND3_X1   g780(.A1(new_n671), .A2(KEYINPUT84), .A3(new_n672), .ZN(new_n1207));
  OAI211_X1 g781(.A(G14), .B(new_n1206), .C1(new_n1207), .C2(new_n674), .ZN(new_n1208));
  NOR2_X1   g782(.A1(G227), .A2(new_n460), .ZN(new_n1209));
  NAND4_X1  g783(.A1(new_n718), .A2(new_n1208), .A3(new_n917), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1205), .A2(new_n1210), .ZN(G308));
  NAND3_X1  g785(.A1(new_n713), .A2(new_n717), .A3(new_n1209), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n1212), .A2(G401), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n1213), .B(new_n917), .C1(new_n992), .C2(new_n993), .ZN(G225));
endmodule


