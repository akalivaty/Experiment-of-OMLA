//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n465), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n473), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n465), .ZN(new_n482));
  INV_X1    g057(.A(G137), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n478), .A2(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n466), .A2(new_n467), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND2_X1  g069(.A1(new_n465), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n471), .B2(new_n473), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n468), .A2(new_n474), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(KEYINPUT4), .C1(new_n486), .C2(new_n495), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n489), .B2(G126), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT71), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G62), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(new_n523), .B1(G75), .B2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(KEYINPUT72), .A3(G62), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n511), .B2(new_n513), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n527), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n526), .A2(new_n534), .ZN(G166));
  INV_X1    g110(.A(new_n531), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  OAI211_X1 g112(.A(G89), .B(new_n521), .C1(new_n529), .C2(new_n530), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(KEYINPUT73), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n538), .B2(new_n540), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n536), .A2(G52), .ZN(new_n546));
  INV_X1    g121(.A(new_n532), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n515), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  XNOR2_X1  g127(.A(KEYINPUT74), .B(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n536), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n547), .A2(G81), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n515), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n521), .A2(G65), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n518), .B2(new_n520), .ZN(new_n570));
  INV_X1    g145(.A(new_n567), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT75), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n568), .A2(G651), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n547), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  OR2_X1    g156(.A1(new_n526), .A2(new_n534), .ZN(G303));
  OAI211_X1 g157(.A(G49), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n583));
  OAI211_X1 g158(.A(G87), .B(new_n521), .C1(new_n529), .C2(new_n530), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n518), .A2(new_n588), .A3(new_n520), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n589), .B2(G651), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n587), .A3(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n586), .A2(new_n593), .ZN(G288));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n518), .B2(new_n520), .ZN(new_n596));
  AND2_X1   g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n514), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g173(.A(G86), .B(new_n521), .C1(new_n529), .C2(new_n530), .ZN(new_n599));
  OAI211_X1 g174(.A(G48), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT77), .ZN(G305));
  NAND2_X1  g177(.A1(new_n536), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT78), .B(G85), .Z(new_n605));
  OAI221_X1 g180(.A(new_n603), .B1(new_n515), .B2(new_n604), .C1(new_n532), .C2(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G301), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n547), .A2(G92), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n531), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(new_n531), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(new_n510), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(KEYINPUT80), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT81), .Z(new_n621));
  AOI21_X1  g196(.A(new_n608), .B1(new_n621), .B2(new_n607), .ZN(G284));
  AOI21_X1  g197(.A(new_n608), .B1(new_n621), .B2(new_n607), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n579), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(G868), .B2(new_n579), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n621), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n621), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n631), .B(new_n632), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g209(.A1(new_n468), .A2(new_n474), .A3(new_n479), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  AOI22_X1  g215(.A1(G123), .A2(new_n489), .B1(new_n487), .B2(G135), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n465), .A2(KEYINPUT83), .A3(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(KEYINPUT83), .B1(new_n465), .B2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT84), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n654), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n667), .A2(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(KEYINPUT85), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(new_n673), .A3(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n667), .B(KEYINPUT17), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n665), .C1(new_n675), .C2(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n669), .A3(new_n664), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n671), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n686), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n688), .B(new_n691), .C1(new_n683), .C2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT88), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n694), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n586), .A2(new_n704), .A3(new_n593), .ZN(new_n705));
  INV_X1    g280(.A(new_n592), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(new_n590), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT91), .B1(new_n707), .B2(new_n585), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT92), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n702), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n702), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n702), .A2(G6), .ZN(new_n720));
  INV_X1    g295(.A(G305), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n702), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n718), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n719), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n713), .A2(KEYINPUT92), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n714), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  OR2_X1    g304(.A1(G95), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT90), .Z(new_n732));
  AOI22_X1  g307(.A1(G119), .A2(new_n489), .B1(new_n487), .B2(G131), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT89), .B(G29), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G25), .B(new_n734), .S(new_n736), .Z(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1986), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n702), .A2(G24), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G290), .B2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n728), .A2(new_n729), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT36), .Z(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT24), .B(G34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n735), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT95), .Z(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G160), .B2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT96), .Z(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G129), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n479), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n762), .B2(G32), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n762), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT25), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n468), .A2(new_n474), .A3(G127), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n465), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n770), .B(new_n773), .C1(G139), .C2(new_n487), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(new_n762), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n765), .A2(new_n767), .B1(G2072), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n753), .B(new_n776), .C1(G2072), .C2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n487), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n489), .A2(G128), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n735), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  INV_X1    g364(.A(G19), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n790), .A2(KEYINPUT93), .A3(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT93), .B1(new_n790), .B2(G16), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n559), .C2(new_n702), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1341), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n736), .A2(G27), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G164), .B2(new_n736), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2078), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n789), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n765), .A2(new_n767), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n702), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n702), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n736), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n736), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT102), .B(KEYINPUT29), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n799), .B1(G1961), .B2(new_n801), .C1(new_n805), .C2(G2090), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n752), .B2(new_n751), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n778), .A2(new_n798), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n702), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n579), .B2(new_n702), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT103), .Z(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(G1956), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(G1956), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n805), .A2(G2090), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT104), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT100), .B1(G16), .B2(G21), .ZN(new_n820));
  NAND2_X1  g395(.A1(G168), .A2(G16), .ZN(new_n821));
  MUX2_X1   g396(.A(KEYINPUT100), .B(new_n820), .S(new_n821), .Z(new_n822));
  INV_X1    g397(.A(G1966), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT31), .B(G11), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(G28), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n762), .B1(new_n827), .B2(G28), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n826), .B1(new_n828), .B2(new_n829), .C1(new_n645), .C2(new_n735), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n801), .B2(G1961), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n824), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n702), .A2(G4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n621), .B2(new_n702), .ZN(new_n835));
  INV_X1    g410(.A(G1348), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n810), .A2(new_n819), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n746), .A2(new_n838), .ZN(G311));
  OR2_X1    g414(.A1(new_n746), .A2(new_n838), .ZN(G150));
  NAND2_X1  g415(.A1(new_n621), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n547), .A2(G93), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT105), .B(G55), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n536), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT106), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT106), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n846), .A2(new_n847), .B1(new_n515), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n558), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n842), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n734), .B(new_n636), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n487), .A2(G142), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n489), .A2(G130), .ZN(new_n860));
  OR2_X1    g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT107), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n508), .B(new_n783), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n761), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n774), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G160), .B(new_n493), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n645), .Z(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n868), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n865), .A2(new_n868), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT40), .Z(G395));
  AND2_X1   g455(.A1(new_n620), .A2(G299), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n611), .B(new_n579), .C1(new_n618), .C2(new_n619), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT41), .B1(new_n881), .B2(new_n883), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n620), .A2(G299), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n849), .B(new_n559), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n629), .B(new_n894), .ZN(new_n895));
  MUX2_X1   g470(.A(new_n885), .B(new_n893), .S(new_n895), .Z(new_n896));
  XOR2_X1   g471(.A(G305), .B(G290), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n709), .B(G166), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n896), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n849), .A2(new_n607), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(G301), .B2(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(G301), .A2(KEYINPUT109), .ZN(new_n913));
  NAND3_X1  g488(.A1(G301), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n912), .A2(new_n913), .A3(G168), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(G168), .B1(KEYINPUT109), .B2(G301), .ZN(new_n916));
  INV_X1    g491(.A(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n911), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n850), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n894), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n891), .A2(new_n892), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n894), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n894), .A3(new_n924), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n884), .A3(new_n919), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n923), .A2(new_n899), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n874), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n899), .B1(new_n923), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n909), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n884), .A2(new_n919), .A3(new_n921), .ZN(new_n933));
  INV_X1    g508(.A(new_n927), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n920), .A2(new_n894), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n934), .A2(new_n925), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n886), .A2(new_n890), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n899), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .A3(new_n874), .A4(new_n929), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n908), .B1(new_n932), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n940), .A2(new_n909), .A3(new_n874), .A4(new_n929), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n908), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n907), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n942), .A2(new_n949), .A3(KEYINPUT112), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(KEYINPUT127), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n783), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT113), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n508), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n484), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n475), .A2(new_n477), .ZN(new_n961));
  OAI211_X1 g536(.A(G40), .B(new_n960), .C1(new_n961), .C2(new_n465), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT114), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n761), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n738), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n734), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n738), .B1(new_n732), .B2(new_n733), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n963), .ZN(new_n973));
  XNOR2_X1  g548(.A(G290), .B(new_n740), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n968), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n478), .A2(new_n979), .A3(new_n484), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n958), .B(G1384), .C1(new_n503), .C2(new_n507), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n717), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n985));
  INV_X1    g560(.A(G2090), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n980), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G166), .B2(new_n978), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT63), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n962), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(new_n752), .A3(new_n988), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n823), .B1(new_n982), .B2(new_n983), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n978), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G168), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n962), .B1(new_n957), .B2(new_n958), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1971), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n980), .B1(new_n981), .B2(new_n987), .ZN(new_n1005));
  AOI211_X1 g580(.A(KEYINPUT50), .B(G1384), .C1(new_n503), .C2(new_n507), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(G2090), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n994), .B(G8), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n990), .A2(KEYINPUT116), .A3(new_n994), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n705), .A2(new_n708), .A3(G1976), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n978), .B1(new_n981), .B2(new_n980), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n601), .A2(new_n1022), .A3(G1981), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n601), .B2(G1981), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1021), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1027), .B(KEYINPUT117), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(KEYINPUT49), .C1(new_n1024), .C2(new_n1023), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1032), .A3(new_n1016), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1020), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1001), .A2(new_n1012), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n984), .A2(new_n989), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT116), .A2(new_n1036), .A3(G8), .A4(new_n994), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n990), .B2(new_n994), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n994), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT119), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n990), .B2(new_n994), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1039), .A2(new_n1045), .A3(new_n1000), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1035), .B1(new_n1046), .B2(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n982), .A2(G2078), .A3(new_n983), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(KEYINPUT53), .ZN(new_n1051));
  INV_X1    g626(.A(G2078), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n959), .A2(new_n1052), .A3(new_n1003), .A4(new_n980), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(G171), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(KEYINPUT53), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(G301), .A4(new_n1049), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(KEYINPUT54), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1056), .A2(KEYINPUT123), .A3(KEYINPUT54), .A4(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n959), .A2(new_n1003), .A3(new_n980), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n575), .B2(new_n578), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n576), .B(KEYINPUT9), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(new_n573), .A3(new_n574), .A4(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n981), .A2(new_n980), .A3(new_n953), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n981), .A2(new_n980), .A3(new_n1078), .A4(new_n953), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n836), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n620), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1074), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1075), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1066), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1084), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1348), .B1(new_n996), .B2(new_n988), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1080), .ZN(new_n1091));
  INV_X1    g666(.A(new_n620), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n1079), .A4(new_n1077), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1074), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1956), .B1(new_n996), .B2(new_n988), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1067), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n982), .A2(new_n983), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1075), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1088), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n982), .A2(G1996), .A3(new_n983), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT58), .B(G1341), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n981), .B2(new_n980), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n559), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT59), .B(new_n559), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1107), .B(new_n1108), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1085), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT54), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1112));
  OAI21_X1  g687(.A(G8), .B1(new_n543), .B2(new_n544), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT122), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(G8), .C1(new_n543), .C2(new_n544), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1966), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1005), .A2(G2084), .A3(new_n1006), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(KEYINPUT51), .C1(new_n999), .C2(new_n1117), .ZN(new_n1121));
  OAI21_X1  g696(.A(G8), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1112), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1064), .A2(new_n1110), .A3(new_n1111), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1012), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1033), .A2(new_n1014), .A3(new_n593), .A4(new_n586), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1031), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1129), .A2(new_n1034), .B1(new_n1131), .B2(new_n1016), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1047), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1121), .A2(KEYINPUT62), .A3(new_n1125), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1012), .A2(new_n1034), .A3(new_n1044), .A4(new_n1042), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT62), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1056), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1137), .A2(new_n1056), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT125), .B1(new_n1141), .B2(new_n1136), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1133), .A2(new_n1134), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1047), .A2(new_n1128), .A3(KEYINPUT124), .A4(new_n1132), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n977), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT48), .Z(new_n1147));
  AND3_X1   g722(.A1(new_n968), .A2(new_n972), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n963), .A2(new_n966), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1150));
  INV_X1    g725(.A(new_n761), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n963), .B1(new_n955), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT47), .Z(new_n1154));
  NOR2_X1   g729(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n968), .A2(new_n970), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n783), .A2(G2067), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT126), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n963), .B1(new_n1158), .B2(KEYINPUT126), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1155), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n952), .B1(new_n1145), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1144), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n977), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1162), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT127), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1163), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(new_n879), .ZN(new_n1173));
  NOR4_X1   g747(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n1173), .A3(new_n1174), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


