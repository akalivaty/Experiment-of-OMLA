//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1326, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  INV_X1    g0005(.A(G50), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G257), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT65), .B(G68), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n205), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n219), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT70), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G107), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n258), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G274), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT71), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AND2_X1   g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n266), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n274), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G244), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n264), .A2(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT74), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n280), .B(new_n286), .C1(new_n281), .C2(new_n283), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n265), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  NAND4_X1  g0089(.A1(KEYINPUT73), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(new_n224), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT73), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n205), .B2(new_n251), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n225), .A2(G1), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(G77), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G20), .A2(G77), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n225), .A2(G33), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n300), .B1(new_n301), .B2(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n293), .A2(new_n224), .A3(new_n290), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n294), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n299), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n265), .A2(G190), .A3(new_n285), .A4(new_n287), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n289), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n285), .A2(new_n287), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n265), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(new_n314), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n280), .B1(new_n207), .B2(new_n283), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n310), .C2(new_n258), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n331), .B2(new_n264), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(G190), .ZN(new_n335));
  INV_X1    g0135(.A(G150), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n301), .A2(new_n304), .B1(new_n336), .B2(new_n303), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n225), .B1(new_n201), .B2(new_n206), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n307), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n298), .A2(G50), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(G50), .B2(new_n294), .C1(new_n295), .C2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT9), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n334), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT10), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n334), .A2(new_n345), .A3(new_n342), .A4(new_n335), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n332), .A2(new_n321), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n341), .B1(new_n332), .B2(G169), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n317), .A2(new_n324), .A3(KEYINPUT76), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n327), .A2(new_n347), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n253), .A2(G33), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT72), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n356), .A2(G232), .A3(G1698), .A4(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n356), .A2(G226), .A3(new_n259), .A4(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n264), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n282), .A2(KEYINPUT77), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n213), .B1(new_n282), .B2(KEYINPUT77), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(new_n279), .B2(new_n271), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n362), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g0168(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT14), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G179), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G68), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT65), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT65), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G68), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT12), .B1(new_n380), .B2(new_n294), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT79), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT12), .A2(G68), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n309), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT79), .B1(new_n385), .B2(new_n294), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n298), .A2(G68), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n295), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT80), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n302), .A2(G50), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n310), .B2(new_n304), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n377), .A2(new_n379), .A3(G20), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT11), .B(new_n307), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n251), .A2(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G77), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n392), .C1(new_n380), .C2(new_n225), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT11), .B1(new_n399), .B2(new_n307), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT80), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n387), .B(new_n402), .C1(new_n295), .C2(new_n389), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n391), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n391), .A2(new_n401), .A3(KEYINPUT81), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n375), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n371), .A2(new_n411), .A3(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n362), .A2(new_n365), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(G190), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(G200), .B1(new_n367), .B2(new_n368), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n410), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n271), .A2(new_n279), .B1(G232), .B2(new_n282), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT82), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n253), .B2(G33), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n251), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n427));
  AND2_X1   g0227(.A1(G226), .A2(G1698), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n254), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT84), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(G223), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1698), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n426), .A2(new_n427), .A3(new_n434), .A4(new_n254), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(G179), .B(new_n424), .C1(new_n438), .C2(new_n267), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n282), .A2(G232), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n268), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n275), .B1(new_n274), .B2(new_n278), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n426), .A2(new_n254), .A3(new_n427), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT84), .A3(new_n428), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n429), .A2(new_n430), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n436), .A4(new_n435), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n447), .B2(new_n264), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n439), .B1(new_n318), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n301), .A2(new_n297), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n296), .A2(new_n450), .B1(new_n309), .B2(new_n301), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT7), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n427), .A2(new_n254), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT82), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n225), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G68), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n426), .A2(new_n254), .A3(new_n427), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n457), .B2(new_n225), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G58), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n202), .B1(new_n214), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(G159), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n303), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(KEYINPUT16), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n307), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g0267(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n252), .A2(new_n254), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n225), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT7), .A2(G20), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n380), .B(new_n472), .C1(new_n258), .C2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n464), .B1(new_n461), .B2(G20), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n451), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n449), .A2(new_n478), .A3(KEYINPUT18), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT85), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n449), .A2(new_n478), .A3(new_n481), .A4(KEYINPUT18), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n449), .A2(new_n478), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT18), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  XOR2_X1   g0286(.A(KEYINPUT86), .B(G190), .Z(new_n487));
  OAI211_X1 g0287(.A(new_n424), .B(new_n487), .C1(new_n438), .C2(new_n267), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G200), .B2(new_n448), .ZN(new_n489));
  INV_X1    g0289(.A(new_n451), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n474), .B1(new_n356), .B2(new_n357), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n452), .B1(new_n470), .B2(new_n225), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n491), .A2(new_n214), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n476), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n307), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n457), .A2(new_n225), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT7), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G68), .A3(new_n455), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT16), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n500), .B(new_n464), .C1(new_n461), .C2(G20), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n496), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n490), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n489), .A2(new_n503), .A3(KEYINPUT17), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT17), .B1(new_n489), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n486), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n353), .A2(new_n423), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G250), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n426), .A2(new_n427), .A3(new_n510), .A4(new_n254), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT92), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G294), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n209), .A2(new_n259), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n426), .A2(new_n515), .A3(new_n254), .A4(new_n427), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n511), .A2(new_n512), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n264), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n277), .A2(G1), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n267), .ZN(new_n524));
  INV_X1    g0324(.A(G264), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT5), .B(G41), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n274), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n519), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n444), .A2(KEYINPUT92), .A3(new_n510), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n526), .B1(new_n533), .B2(new_n264), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n534), .B2(new_n529), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n426), .A2(new_n427), .A3(new_n225), .A4(new_n254), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT22), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n538), .A2(KEYINPUT22), .A3(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n356), .A2(new_n357), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n225), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n262), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n545), .A2(new_n546), .B1(new_n548), .B2(new_n225), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n543), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n307), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n309), .A2(new_n262), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT25), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n269), .A2(G33), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n291), .A2(new_n293), .A3(new_n294), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n554), .B1(G107), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT94), .B1(new_n536), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n552), .A2(new_n558), .ZN(new_n561));
  INV_X1    g0361(.A(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n534), .A2(new_n562), .A3(new_n529), .ZN(new_n563));
  INV_X1    g0363(.A(new_n530), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(G200), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT94), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n530), .A2(G169), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n534), .A2(G179), .A3(new_n529), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT93), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n559), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n294), .A2(G97), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n557), .B2(G97), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n579), .A2(new_n208), .A3(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n582), .A2(new_n225), .B1(new_n310), .B2(new_n303), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n472), .B1(new_n258), .B2(new_n474), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n262), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n578), .B1(new_n586), .B2(new_n307), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n509), .B2(new_n259), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n356), .A2(new_n357), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G283), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n281), .A2(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n426), .A2(new_n427), .A3(new_n592), .A4(new_n254), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n264), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n523), .A2(G257), .A3(new_n267), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n529), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n529), .A3(new_n598), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(G190), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n599), .A2(new_n598), .A3(new_n529), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n600), .ZN(new_n606));
  AOI21_X1  g0406(.A(G200), .B1(new_n606), .B2(new_n597), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n587), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n318), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n491), .A2(new_n262), .A3(new_n492), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n307), .B1(new_n610), .B2(new_n583), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n577), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n321), .A3(new_n597), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G303), .B1(new_n256), .B2(new_n257), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n525), .A2(G1698), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G257), .B2(G1698), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n444), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n267), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G270), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n529), .B1(new_n524), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT21), .B(G169), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G303), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n356), .B2(new_n357), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n457), .A2(new_n618), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n264), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(G179), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n557), .A2(G116), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT20), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(KEYINPUT91), .ZN(new_n634));
  AOI21_X1  g0434(.A(G20), .B1(G33), .B2(G283), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n251), .A2(G97), .ZN(new_n636));
  INV_X1    g0436(.A(G116), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n635), .A2(new_n636), .B1(G20), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n307), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n633), .A2(KEYINPUT91), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n309), .A2(KEYINPUT90), .A3(new_n637), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n294), .B2(G116), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n307), .A2(KEYINPUT91), .A3(new_n638), .A4(new_n633), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n632), .A2(new_n642), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n631), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n628), .A2(new_n629), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G200), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n556), .B2(new_n637), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n634), .B(new_n640), .C1(new_n307), .C2(new_n638), .ZN(new_n653));
  INV_X1    g0453(.A(new_n647), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n655), .C1(new_n487), .C2(new_n650), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n318), .B1(new_n628), .B2(new_n629), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n648), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT21), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n649), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT19), .ZN(new_n662));
  NOR2_X1   g0462(.A1(G97), .A2(G107), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n538), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n360), .A2(new_n225), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n304), .A2(KEYINPUT19), .A3(new_n208), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n537), .B2(new_n376), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n496), .B1(new_n668), .B2(KEYINPUT88), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n397), .A2(new_n662), .A3(G97), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n663), .A2(new_n538), .B1(new_n360), .B2(new_n225), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n662), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n672), .B(new_n673), .C1(new_n376), .C2(new_n537), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n669), .A2(new_n674), .B1(new_n309), .B2(new_n305), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n267), .A2(G274), .A3(new_n520), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n269), .A2(G45), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n267), .A2(G250), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n281), .A2(G1698), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(G238), .B2(G1698), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n547), .B1(new_n457), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(new_n264), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G190), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT89), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n556), .A2(new_n538), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n264), .ZN(new_n687));
  INV_X1    g0487(.A(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n686), .B1(new_n689), .B2(G200), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT89), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n683), .A2(new_n691), .A3(G190), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n675), .A2(new_n685), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n307), .A3(new_n674), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n305), .A2(new_n309), .ZN(new_n696));
  INV_X1    g0496(.A(new_n305), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n557), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AOI211_X1 g0499(.A(G179), .B(new_n679), .C1(new_n264), .C2(new_n682), .ZN(new_n700));
  AOI21_X1  g0500(.A(G169), .B1(new_n687), .B2(new_n688), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n615), .A2(new_n661), .A3(new_n704), .ZN(new_n705));
  AND4_X1   g0505(.A1(new_n508), .A2(new_n568), .A3(new_n575), .A4(new_n705), .ZN(G372));
  AND3_X1   g0506(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n707), .A2(new_n321), .B1(new_n611), .B2(new_n577), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n609), .A3(new_n693), .A4(new_n703), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(KEYINPUT26), .B1(new_n699), .B2(new_n702), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT26), .ZN(new_n711));
  INV_X1    g0511(.A(new_n614), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n675), .A2(new_n690), .A3(new_n684), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n703), .A2(new_n713), .A3(KEYINPUT95), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT95), .B1(new_n703), .B2(new_n713), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n711), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n571), .A2(new_n559), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n649), .B2(new_n660), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n655), .B1(new_n624), .B2(new_n630), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT21), .B1(new_n657), .B2(new_n648), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT96), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n718), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n608), .A2(new_n614), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n703), .A2(new_n713), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n703), .A2(new_n713), .A3(KEYINPUT95), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n568), .A2(new_n724), .A3(new_n725), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n717), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n508), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n485), .A2(new_n479), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n422), .A2(new_n735), .B1(new_n375), .B2(new_n409), .ZN(new_n736));
  INV_X1    g0536(.A(new_n506), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n350), .B1(new_n738), .B2(new_n347), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(new_n739), .ZN(G369));
  NOR2_X1   g0540(.A1(new_n720), .A2(new_n723), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n269), .A2(new_n225), .A3(G13), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT27), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT27), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(G213), .ZN(new_n745));
  INV_X1    g0545(.A(G343), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n655), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n741), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n661), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT97), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n536), .A2(KEYINPUT94), .A3(new_n559), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n566), .B1(new_n561), .B2(new_n565), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n575), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n561), .A2(new_n748), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n559), .A2(new_n747), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n568), .A2(KEYINPUT97), .A3(new_n575), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n575), .A2(new_n748), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n752), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n721), .A2(new_n722), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n747), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n758), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n571), .A2(new_n559), .A3(new_n748), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n764), .A2(new_n769), .ZN(G399));
  INV_X1    g0570(.A(new_n221), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT98), .B1(new_n771), .B2(G41), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n771), .A2(KEYINPUT98), .A3(G41), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n663), .A2(new_n538), .A3(new_n637), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n775), .A2(new_n269), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n229), .B2(new_n775), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  AOI21_X1  g0579(.A(new_n747), .B1(new_n717), .B2(new_n731), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(KEYINPUT29), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n703), .B1(new_n709), .B2(KEYINPUT26), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n730), .A2(new_n712), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(KEYINPUT26), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n575), .A2(new_n765), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n785), .A2(new_n568), .A3(new_n725), .A4(new_n730), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n747), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n781), .B1(KEYINPUT29), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G330), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n705), .A2(new_n568), .A3(new_n575), .A4(new_n748), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT30), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n529), .B(G179), .C1(new_n524), .C2(new_n622), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n621), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n793), .A2(new_n597), .A3(new_n606), .A4(new_n683), .ZN(new_n794));
  INV_X1    g0594(.A(new_n534), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n689), .A2(new_n621), .A3(new_n792), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n707), .A2(new_n797), .A3(KEYINPUT30), .A4(new_n534), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n683), .A2(G179), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n530), .A2(new_n603), .A3(new_n650), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  AND3_X1   g0601(.A1(new_n801), .A2(KEYINPUT31), .A3(new_n747), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT31), .B1(new_n801), .B2(new_n747), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n789), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n779), .B1(new_n806), .B2(G1), .ZN(G364));
  INV_X1    g0607(.A(new_n752), .ZN(new_n808));
  INV_X1    g0608(.A(G13), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n269), .B1(new_n810), .B2(G45), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n775), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G330), .B2(new_n751), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n224), .B1(G20), .B2(new_n318), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n225), .A2(new_n321), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G200), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n487), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT100), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G50), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n225), .A2(G179), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G190), .A2(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n463), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT32), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n829), .A2(new_n562), .A3(G200), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n258), .B1(new_n262), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n819), .A2(new_n830), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n840), .B2(G77), .ZN(new_n841));
  INV_X1    g0641(.A(new_n819), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n487), .A2(new_n842), .A3(G200), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n829), .A2(G190), .A3(G200), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n844), .A2(new_n460), .B1(new_n538), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n820), .A2(G190), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n562), .A2(G179), .A3(G200), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n225), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n848), .A2(new_n376), .B1(new_n208), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n828), .A2(new_n833), .A3(new_n841), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT101), .B(G326), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n827), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(KEYINPUT33), .A2(G317), .ZN(new_n856));
  AND2_X1   g0656(.A1(KEYINPUT33), .A2(G317), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G294), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n850), .ZN(new_n860));
  INV_X1    g0660(.A(new_n834), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(G283), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n819), .A2(G311), .A3(new_n830), .ZN(new_n863));
  INV_X1    g0663(.A(new_n831), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n863), .B(new_n258), .C1(G329), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n845), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n843), .A2(G322), .B1(new_n866), .B2(G303), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n855), .A2(new_n862), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n818), .B1(new_n853), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(G13), .A2(G33), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(G20), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n817), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n258), .A2(G355), .A3(new_n221), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n249), .A2(G45), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n444), .A2(new_n771), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(G45), .B2(new_n228), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n874), .B1(G116), .B2(new_n221), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n816), .B(new_n869), .C1(new_n873), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n872), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n751), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n815), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G396));
  NOR2_X1   g0683(.A1(new_n324), .A2(new_n747), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n323), .A2(new_n747), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n316), .A2(new_n314), .A3(new_n315), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n333), .B1(new_n320), .B2(new_n265), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n324), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n780), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n780), .A2(new_n889), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n805), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n813), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n805), .A3(new_n891), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n817), .A2(new_n870), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n816), .B1(new_n310), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n861), .A2(G87), .ZN(new_n898));
  INV_X1    g0698(.A(G283), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n898), .B1(new_n848), .B2(new_n899), .C1(new_n844), .C2(new_n859), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n258), .B1(G311), .B2(new_n864), .ZN(new_n901));
  INV_X1    g0701(.A(new_n850), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n902), .A2(G97), .B1(new_n866), .B2(G107), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n901), .B(new_n903), .C1(new_n637), .C2(new_n839), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n900), .B(new_n904), .C1(G303), .C2(new_n827), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n843), .A2(G143), .B1(new_n847), .B2(G150), .ZN(new_n906));
  INV_X1    g0706(.A(G137), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n906), .B1(new_n463), .B2(new_n839), .C1(new_n826), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT34), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n850), .A2(new_n460), .B1(new_n834), .B2(new_n376), .ZN(new_n910));
  INV_X1    g0710(.A(G132), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n444), .B1(new_n911), .B2(new_n831), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n910), .B(new_n912), .C1(G50), .C2(new_n866), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n905), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n897), .B1(new_n818), .B2(new_n914), .C1(new_n889), .C2(new_n871), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n895), .A2(new_n915), .ZN(G384));
  NOR2_X1   g0716(.A1(new_n810), .A2(new_n269), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n485), .A2(new_n479), .A3(new_n745), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n469), .B1(new_n499), .B2(new_n476), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n451), .B1(new_n467), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT104), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(new_n451), .C1(new_n467), .C2(new_n921), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n439), .B(new_n745), .C1(new_n318), .C2(new_n448), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n489), .A2(new_n503), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n920), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n483), .A2(new_n928), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  INV_X1    g0731(.A(new_n745), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n478), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n930), .A2(new_n931), .A3(new_n920), .A4(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n483), .A2(new_n928), .A3(new_n933), .A4(new_n920), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n929), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n923), .A2(new_n932), .A3(new_n925), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n486), .B2(new_n506), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n919), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n927), .A2(new_n928), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n938), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n507), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT38), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n940), .A2(new_n948), .A3(KEYINPUT106), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT106), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n919), .C1(new_n937), .C2(new_n939), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n735), .A2(new_n748), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n891), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n420), .B1(new_n412), .B2(new_n417), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n409), .B(new_n747), .C1(new_n955), .C2(new_n375), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n409), .A2(new_n747), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n410), .A2(new_n422), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n949), .A2(KEYINPUT39), .A3(new_n951), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n483), .A2(new_n928), .A3(new_n933), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n934), .A2(new_n936), .B1(KEYINPUT37), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n933), .B1(new_n506), .B2(new_n734), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n919), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n948), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n961), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n375), .A2(new_n409), .A3(new_n748), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n918), .B1(new_n952), .B2(new_n960), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n784), .A2(new_n786), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(KEYINPUT29), .A3(new_n748), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n508), .C1(KEYINPUT29), .C2(new_n780), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n739), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n970), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n965), .A2(new_n948), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n888), .A2(new_n324), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n953), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n790), .B2(new_n804), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(KEYINPUT40), .A3(new_n959), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n976), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n980), .A2(KEYINPUT40), .A3(new_n959), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n965), .A2(new_n948), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(KEYINPUT107), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n949), .A2(new_n951), .A3(new_n959), .A4(new_n980), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT40), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n508), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n790), .B2(new_n804), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n789), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n990), .B2(new_n992), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n917), .B1(new_n975), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n975), .B2(new_n994), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n310), .B(new_n228), .C1(new_n380), .C2(G58), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n206), .A2(G68), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT103), .Z(new_n999));
  OAI211_X1 g0799(.A(G1), .B(new_n809), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n582), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT35), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT35), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1002), .A2(G116), .A3(new_n227), .A4(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n996), .A2(new_n1000), .A3(new_n1006), .ZN(G367));
  NAND2_X1  g0807(.A1(new_n761), .A2(new_n763), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n808), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n725), .B1(new_n587), .B2(new_n748), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n712), .A2(new_n747), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT108), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n764), .A2(new_n1015), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n675), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n747), .B1(new_n1018), .B2(new_n686), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n730), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n703), .B2(new_n1019), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n1017), .A2(KEYINPUT43), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n767), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n1012), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT42), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n614), .B1(new_n1010), .B2(new_n575), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1024), .A2(KEYINPUT42), .B1(new_n748), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1025), .A2(new_n1027), .B1(KEYINPUT43), .B2(new_n1021), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1017), .B1(KEYINPUT43), .B2(new_n1021), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1022), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1028), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n775), .B(KEYINPUT41), .Z(new_n1033));
  NAND3_X1  g0833(.A1(new_n767), .A2(new_n768), .A3(new_n1012), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT45), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT44), .B1(new_n769), .B2(new_n1013), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n769), .A2(new_n1013), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT44), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1036), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n764), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n762), .B(new_n766), .C1(new_n758), .C2(new_n760), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n808), .B1(new_n1043), .B2(new_n1023), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n752), .B(new_n767), .C1(new_n1008), .C2(new_n766), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n806), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT109), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1038), .B(new_n1039), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n1009), .A3(new_n1036), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT109), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n806), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1042), .A2(new_n1048), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n1053), .B2(new_n806), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1032), .B1(new_n1054), .B2(new_n812), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n834), .A2(new_n208), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n844), .A2(new_n625), .B1(new_n848), .B2(new_n859), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G107), .C2(new_n902), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n866), .A2(G116), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT46), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT111), .B(G317), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n444), .B(new_n1061), .C1(new_n864), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n827), .A2(G311), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n840), .A2(G283), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1058), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n827), .A2(G143), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n844), .A2(new_n336), .B1(new_n460), .B2(new_n845), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G159), .B2(new_n847), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n840), .A2(G50), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n356), .A2(new_n357), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n850), .A2(new_n376), .B1(new_n834), .B2(new_n310), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G137), .C2(new_n864), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT47), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT47), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n817), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n241), .A2(new_n876), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n873), .B1(new_n221), .B2(new_n305), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n813), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT110), .Z(new_n1082));
  OAI211_X1 g0882(.A(new_n1078), .B(new_n1082), .C1(new_n1021), .C2(new_n880), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1055), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT112), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G387));
  NAND3_X1  g0886(.A1(new_n258), .A2(new_n221), .A3(new_n776), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n876), .B1(new_n236), .B2(new_n277), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n301), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1089), .A2(KEYINPUT50), .A3(new_n206), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT50), .B1(new_n1089), .B2(new_n206), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n277), .B1(new_n376), .B2(new_n310), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n776), .B2(KEYINPUT113), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(KEYINPUT113), .B2(new_n776), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1087), .B1(G107), .B2(new_n221), .C1(new_n1088), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n873), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n813), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n843), .A2(new_n1062), .B1(new_n847), .B2(G311), .ZN(new_n1100));
  INV_X1    g0900(.A(G322), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1100), .B1(new_n625), .B2(new_n839), .C1(new_n826), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT48), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n902), .A2(G283), .B1(new_n866), .B2(G294), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT49), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n444), .B1(new_n854), .B2(new_n864), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n637), .B2(new_n834), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n848), .A2(new_n301), .B1(new_n208), .B2(new_n834), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n836), .A2(new_n376), .B1(new_n831), .B2(new_n336), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n457), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n845), .A2(new_n310), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n843), .B2(G50), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(new_n305), .C2(new_n850), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G159), .B2(new_n827), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1099), .B1(new_n1122), .B2(new_n817), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT114), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n1008), .C2(new_n880), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n813), .B(new_n1098), .C1(new_n1126), .C2(new_n818), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1008), .A2(new_n880), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT114), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1125), .A2(new_n1129), .B1(new_n1046), .B2(new_n812), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1044), .B(new_n1045), .C1(new_n788), .C2(new_n805), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1047), .A2(new_n775), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(G393));
  INV_X1    g0933(.A(new_n1050), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1009), .B1(new_n1049), .B2(new_n1036), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1047), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n1053), .A3(new_n775), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1042), .A2(new_n812), .A3(new_n1050), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n246), .A2(new_n876), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n873), .B1(new_n208), .B2(new_n221), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n813), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n827), .A2(G317), .B1(G311), .B2(new_n843), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT52), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1071), .B1(new_n859), .B2(new_n836), .C1(new_n1101), .C2(new_n831), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n847), .A2(G303), .B1(new_n861), .B2(G107), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n637), .B2(new_n850), .C1(new_n899), .C2(new_n845), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n826), .A2(new_n336), .B1(new_n463), .B2(new_n844), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT51), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n840), .A2(new_n1089), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G77), .A2(new_n902), .B1(new_n847), .B2(G50), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1150), .A2(new_n444), .A3(new_n898), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G143), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n845), .A2(new_n214), .B1(new_n831), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT115), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1149), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT116), .Z(new_n1158));
  AOI21_X1  g0958(.A(new_n1141), .B1(new_n1158), .B2(new_n817), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n880), .B2(new_n1012), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1138), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1137), .A2(new_n1161), .ZN(G390));
  AOI21_X1  g0962(.A(new_n884), .B1(new_n780), .B2(new_n889), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n956), .A2(new_n958), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n969), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n961), .A3(new_n967), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n969), .B(KEYINPUT117), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n884), .B1(new_n787), .B2(new_n978), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n984), .B(new_n1167), .C1(new_n1168), .C2(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n805), .A2(new_n959), .A3(new_n889), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1166), .A2(new_n1171), .A3(new_n1169), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n508), .A2(new_n805), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n973), .A2(new_n739), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n661), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n704), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n725), .A2(new_n1178), .A3(new_n1179), .A4(new_n748), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n756), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n803), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n801), .A2(KEYINPUT31), .A3(new_n747), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G330), .B(new_n889), .C1(new_n1181), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1164), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT118), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1164), .A3(KEYINPUT118), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1188), .A2(new_n1171), .A3(new_n1168), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1171), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n954), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1177), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1175), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1173), .A2(new_n1174), .A3(new_n1193), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n775), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1173), .A2(new_n812), .A3(new_n1174), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT120), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n896), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n813), .B1(new_n1089), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n827), .A2(G283), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n844), .A2(new_n637), .B1(new_n310), .B2(new_n850), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G107), .B2(new_n847), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n840), .A2(G97), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n834), .A2(new_n376), .B1(new_n845), .B2(new_n538), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n258), .B(new_n1206), .C1(G294), .C2(new_n864), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n258), .B1(new_n206), .B2(new_n834), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n845), .A2(new_n336), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT53), .ZN(new_n1212));
  INV_X1    g1012(.A(G128), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1210), .B(new_n1212), .C1(new_n1213), .C2(new_n826), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n843), .A2(G132), .B1(new_n847), .B2(G137), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n902), .A2(G159), .B1(G125), .B2(new_n864), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT54), .B(G143), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1216), .C1(new_n839), .C2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1208), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1201), .B1(new_n1219), .B2(new_n817), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n961), .A2(new_n967), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n871), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1198), .A2(new_n1199), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1199), .B1(new_n1198), .B2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1197), .B1(new_n1223), .B2(new_n1224), .ZN(G378));
  NAND2_X1  g1025(.A1(new_n347), .A2(new_n351), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n341), .A2(new_n932), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1226), .B(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1228), .B(new_n1229), .ZN(new_n1230));
  AND4_X1   g1030(.A1(G330), .A2(new_n986), .A3(new_n989), .A4(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n789), .B1(new_n982), .B2(new_n985), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1232), .B2(new_n989), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n970), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1230), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n983), .A2(KEYINPUT107), .A3(new_n984), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT107), .B1(new_n983), .B2(new_n984), .ZN(new_n1237));
  OAI21_X1  g1037(.A(G330), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n989), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n918), .B1(new_n960), .B2(new_n952), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n969), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n1221), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1232), .A2(new_n989), .A3(new_n1230), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1234), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n812), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1235), .A2(new_n870), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n813), .B1(G50), .B2(new_n1200), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n848), .A2(new_n911), .B1(new_n836), .B2(new_n907), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT122), .Z(new_n1251));
  NAND2_X1  g1051(.A1(new_n827), .A2(G125), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n850), .A2(new_n336), .B1(new_n845), .B2(new_n1217), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G128), .B2(new_n843), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(KEYINPUT59), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT59), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n861), .A2(G159), .ZN(new_n1258));
  AOI211_X1 g1058(.A(G33), .B(G41), .C1(new_n864), .C2(G124), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1118), .B1(G68), .B2(new_n902), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n460), .B2(new_n834), .C1(new_n262), .C2(new_n844), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n276), .B1(new_n831), .B2(new_n899), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1262), .A2(new_n444), .A3(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n848), .A2(new_n208), .B1(new_n305), .B2(new_n836), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT121), .Z(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n637), .C2(new_n826), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT58), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n276), .B1(new_n457), .B2(new_n251), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n206), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1260), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1249), .B1(new_n1273), .B2(new_n817), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1248), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1247), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1177), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1196), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n775), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1234), .B2(new_n1245), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n1278), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1276), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(G375));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n811), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1164), .A2(new_n870), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n813), .B1(G68), .B2(new_n1200), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n843), .A2(G283), .B1(new_n866), .B2(G97), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n637), .B2(new_n848), .C1(new_n826), .C2(new_n859), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n258), .B1(G303), .B2(new_n864), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n902), .A2(new_n697), .B1(new_n861), .B2(G77), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1293), .B(new_n1294), .C1(new_n262), .C2(new_n839), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n826), .A2(new_n911), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n848), .A2(new_n1217), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n902), .A2(G50), .B1(new_n866), .B2(G159), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n843), .A2(G137), .B1(new_n861), .B2(G58), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n836), .A2(new_n336), .B1(new_n831), .B2(new_n1213), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n457), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n1292), .A2(new_n1295), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1290), .B1(new_n1303), .B2(new_n817), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1289), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1287), .B1(new_n1288), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1163), .B1(new_n1171), .B2(new_n1186), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1185), .A2(new_n1164), .A3(KEYINPUT118), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT118), .B1(new_n1185), .B2(new_n1164), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(KEYINPUT123), .B(new_n1305), .C1(new_n1313), .C2(new_n811), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1033), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1190), .A2(new_n1177), .A3(new_n1192), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1194), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(G381));
  AND2_X1   g1119(.A1(new_n1198), .A2(new_n1222), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1197), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1130), .A2(new_n1132), .A3(new_n882), .ZN(new_n1323));
  NOR4_X1   g1123(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1085), .A2(new_n1285), .A3(new_n1322), .A4(new_n1324), .ZN(G407));
  NAND3_X1  g1125(.A1(new_n1285), .A2(new_n746), .A3(new_n1322), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G407), .A2(G213), .A3(new_n1326), .ZN(G409));
  AND2_X1   g1127(.A1(new_n746), .A2(G213), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n1246), .A2(new_n812), .B1(new_n1248), .B2(new_n1274), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1240), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1243), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1278), .B(KEYINPUT57), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n775), .ZN(new_n1333));
  OAI211_X1 g1133(.A(G378), .B(new_n1329), .C1(new_n1333), .C2(new_n1279), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1246), .A2(new_n1316), .A3(new_n1278), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1247), .A3(new_n1275), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1322), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1328), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT60), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1317), .B1(new_n1193), .B2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1190), .A2(new_n1177), .A3(KEYINPUT60), .A4(new_n1192), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1341), .A2(new_n775), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1343), .A2(new_n1315), .A3(G384), .ZN(new_n1344));
  AOI21_X1  g1144(.A(G384), .B1(new_n1343), .B2(new_n1315), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT124), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(G384), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1307), .A2(new_n1314), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1341), .A2(new_n775), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT60), .B1(new_n1313), .B2(new_n1177), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1350), .B1(new_n1351), .B2(new_n1317), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1348), .B1(new_n1349), .B2(new_n1352), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1343), .A2(new_n1315), .A3(G384), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT124), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  OR2_X1    g1155(.A1(new_n1347), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1338), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT63), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1328), .A2(G2897), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1360), .B1(new_n1347), .B2(new_n1355), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1362), .A2(G2897), .A3(new_n1328), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1364));
  OR2_X1    g1164(.A1(new_n1338), .A2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1356), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n882), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(KEYINPUT112), .B1(new_n1368), .B2(new_n1323), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(G390), .A2(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1323), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1371), .A2(new_n1367), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1372), .B1(new_n1137), .B2(new_n1161), .ZN(new_n1373));
  OAI211_X1 g1173(.A(new_n1055), .B(new_n1083), .C1(new_n1370), .C2(new_n1373), .ZN(new_n1374));
  OAI21_X1  g1174(.A(G390), .B1(new_n1371), .B2(new_n1367), .ZN(new_n1375));
  OAI211_X1 g1175(.A(new_n1137), .B(new_n1161), .C1(new_n1372), .C2(KEYINPUT112), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1084), .A2(new_n1375), .A3(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1374), .A2(new_n1377), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1378), .A2(KEYINPUT61), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1359), .A2(new_n1365), .A3(new_n1366), .A4(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT62), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1338), .A2(new_n1381), .A3(new_n1356), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1383), .B1(new_n1338), .B2(new_n1364), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1381), .B1(new_n1338), .B2(new_n1356), .ZN(new_n1385));
  NOR3_X1   g1185(.A1(new_n1382), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1378), .ZN(new_n1387));
  OAI21_X1  g1187(.A(new_n1380), .B1(new_n1386), .B2(new_n1387), .ZN(G405));
  INV_X1    g1188(.A(KEYINPUT126), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1334), .ZN(new_n1390));
  AOI22_X1  g1190(.A1(new_n1234), .A2(new_n1245), .B1(new_n1277), .B2(new_n1196), .ZN(new_n1391));
  OAI211_X1 g1191(.A(new_n1332), .B(new_n775), .C1(new_n1391), .C2(KEYINPUT57), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1321), .B1(new_n1392), .B2(new_n1329), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1389), .B1(new_n1390), .B2(new_n1393), .ZN(new_n1394));
  OAI211_X1 g1194(.A(KEYINPUT126), .B(new_n1334), .C1(new_n1285), .C2(new_n1321), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1394), .A2(new_n1356), .A3(new_n1395), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1374), .A2(new_n1377), .A3(KEYINPUT127), .ZN(new_n1397));
  OAI211_X1 g1197(.A(new_n1334), .B(new_n1362), .C1(new_n1285), .C2(new_n1321), .ZN(new_n1398));
  AND2_X1   g1198(.A1(new_n1397), .A2(new_n1398), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1396), .A2(new_n1399), .ZN(new_n1400));
  NOR2_X1   g1200(.A1(new_n1387), .A2(KEYINPUT127), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1400), .A2(new_n1401), .ZN(new_n1402));
  OAI211_X1 g1202(.A(new_n1396), .B(new_n1399), .C1(KEYINPUT127), .C2(new_n1387), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1402), .A2(new_n1403), .ZN(G402));
endmodule


