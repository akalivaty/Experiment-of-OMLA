

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n730), .ZN(n714) );
  BUF_X1 U549 ( .A(n604), .Z(n605) );
  XNOR2_X1 U550 ( .A(KEYINPUT65), .B(G2104), .ZN(n525) );
  NAND2_X2 U551 ( .A1(n685), .A2(n772), .ZN(n730) );
  XNOR2_X1 U552 ( .A(n527), .B(n526), .ZN(n604) );
  INV_X1 U553 ( .A(KEYINPUT67), .ZN(n526) );
  NOR2_X1 U554 ( .A1(n525), .A2(G2105), .ZN(n527) );
  NOR2_X1 U555 ( .A1(n697), .A2(n912), .ZN(n692) );
  INV_X1 U556 ( .A(n917), .ZN(n749) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n769) );
  NOR2_X1 U558 ( .A1(n541), .A2(n540), .ZN(G160) );
  AND2_X1 U559 ( .A1(n809), .A2(n800), .ZN(n513) );
  NAND2_X1 U560 ( .A1(G286), .A2(G8), .ZN(n514) );
  OR2_X1 U561 ( .A1(n764), .A2(n753), .ZN(n515) );
  NOR2_X1 U562 ( .A1(n764), .A2(n749), .ZN(n516) );
  NAND2_X1 U563 ( .A1(n730), .A2(G1341), .ZN(n688) );
  INV_X1 U564 ( .A(KEYINPUT95), .ZN(n700) );
  XNOR2_X1 U565 ( .A(n700), .B(KEYINPUT27), .ZN(n701) );
  XNOR2_X1 U566 ( .A(n702), .B(n701), .ZN(n704) );
  AND2_X1 U567 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U568 ( .A(n739), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U569 ( .A1(n927), .A2(n515), .ZN(n754) );
  XNOR2_X1 U570 ( .A(n517), .B(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U571 ( .A(n519), .B(n518), .ZN(n534) );
  INV_X1 U572 ( .A(KEYINPUT66), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n513), .A2(n801), .ZN(n802) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n646) );
  OR2_X1 U575 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U576 ( .A1(G651), .A2(n642), .ZN(n654) );
  XNOR2_X1 U577 ( .A(KEYINPUT23), .B(n533), .ZN(n541) );
  NOR2_X1 U578 ( .A1(n532), .A2(n531), .ZN(G164) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  INV_X1 U580 ( .A(KEYINPUT68), .ZN(n517) );
  INV_X1 U581 ( .A(n534), .ZN(n520) );
  INV_X1 U582 ( .A(n520), .ZN(n865) );
  NAND2_X1 U583 ( .A1(G138), .A2(n865), .ZN(n522) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n868) );
  NAND2_X1 U585 ( .A1(n868), .A2(G114), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n525), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U588 ( .A(n524), .B(n523), .ZN(n869) );
  NAND2_X1 U589 ( .A1(G126), .A2(n869), .ZN(n530) );
  NAND2_X1 U590 ( .A1(G102), .A2(n604), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT88), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U593 ( .A1(n604), .A2(G101), .ZN(n533) );
  NAND2_X1 U594 ( .A1(G137), .A2(n534), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G113), .A2(n868), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U597 ( .A(n537), .B(KEYINPUT69), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G125), .A2(n869), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  INV_X1 U603 ( .A(G108), .ZN(G238) );
  NAND2_X1 U604 ( .A1(G90), .A2(n646), .ZN(n544) );
  INV_X1 U605 ( .A(G651), .ZN(n547) );
  XOR2_X1 U606 ( .A(G543), .B(KEYINPUT0), .Z(n542) );
  XNOR2_X1 U607 ( .A(KEYINPUT70), .B(n542), .ZN(n642) );
  NOR2_X1 U608 ( .A1(n547), .A2(n642), .ZN(n649) );
  NAND2_X1 U609 ( .A1(G77), .A2(n649), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT9), .B(n545), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n654), .A2(G52), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT72), .ZN(n550) );
  NOR2_X1 U614 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n548), .Z(n645) );
  NAND2_X1 U616 ( .A1(G64), .A2(n645), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT73), .B(n551), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(G301) );
  NAND2_X1 U620 ( .A1(n646), .A2(G89), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G76), .A2(n649), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT5), .B(n557), .ZN(n565) );
  XNOR2_X1 U625 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n645), .A2(G63), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n558), .B(KEYINPUT76), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G51), .A2(n654), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(KEYINPUT6), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(n566), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n819) );
  NAND2_X1 U638 ( .A1(n819), .A2(G567), .ZN(n568) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  XOR2_X1 U640 ( .A(G860), .B(KEYINPUT74), .Z(n598) );
  NAND2_X1 U641 ( .A1(G56), .A2(n645), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n569), .Z(n575) );
  NAND2_X1 U643 ( .A1(n646), .A2(G81), .ZN(n570) );
  XNOR2_X1 U644 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U645 ( .A1(G68), .A2(n649), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n654), .A2(G43), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n932) );
  OR2_X1 U651 ( .A1(n598), .A2(n932), .ZN(G153) );
  NAND2_X1 U652 ( .A1(G54), .A2(n654), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G79), .A2(n649), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G66), .A2(n645), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G92), .A2(n646), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT15), .ZN(n912) );
  INV_X1 U660 ( .A(n912), .ZN(n616) );
  NOR2_X1 U661 ( .A1(n616), .A2(G868), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT75), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G65), .A2(n645), .ZN(n589) );
  NAND2_X1 U666 ( .A1(G53), .A2(n654), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G91), .A2(n646), .ZN(n591) );
  NAND2_X1 U669 ( .A1(G78), .A2(n649), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n708) );
  INV_X1 U672 ( .A(n708), .ZN(G299) );
  XNOR2_X1 U673 ( .A(KEYINPUT79), .B(G868), .ZN(n594) );
  NOR2_X1 U674 ( .A1(G286), .A2(n594), .ZN(n597) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n595), .B(KEYINPUT80), .ZN(n596) );
  NOR2_X1 U677 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n599), .A2(n616), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n932), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G868), .A2(n616), .ZN(n601) );
  NOR2_X1 U683 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U684 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G111), .A2(n868), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G99), .A2(n605), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G123), .A2(n869), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G135), .A2(n865), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT81), .B(n611), .Z(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n975) );
  XNOR2_X1 U694 ( .A(G2096), .B(n975), .ZN(n615) );
  INV_X1 U695 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U697 ( .A1(n616), .A2(G559), .ZN(n664) );
  XNOR2_X1 U698 ( .A(n932), .B(n664), .ZN(n617) );
  NOR2_X1 U699 ( .A1(G860), .A2(n617), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G67), .A2(n645), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G55), .A2(n654), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G93), .A2(n646), .ZN(n621) );
  NAND2_X1 U704 ( .A1(G80), .A2(n649), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n667) );
  XNOR2_X1 U707 ( .A(n667), .B(KEYINPUT82), .ZN(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U709 ( .A1(n654), .A2(G47), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n645), .A2(G60), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U712 ( .A(KEYINPUT71), .B(n628), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G85), .A2(n646), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G72), .A2(n649), .ZN(n629) );
  AND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G88), .A2(n646), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G75), .A2(n649), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G62), .A2(n645), .ZN(n636) );
  NAND2_X1 U721 ( .A1(G50), .A2(n654), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U723 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G49), .A2(n654), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U727 ( .A1(n645), .A2(n641), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G87), .A2(n642), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G61), .A2(n645), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G86), .A2(n646), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n653) );
  NAND2_X1 U733 ( .A1(G73), .A2(n649), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n650), .B(KEYINPUT83), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n651), .B(KEYINPUT2), .ZN(n652) );
  NOR2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n654), .A2(G48), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(G305) );
  XNOR2_X1 U739 ( .A(G290), .B(n932), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n658) );
  XNOR2_X1 U741 ( .A(n708), .B(G166), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n659), .B(G288), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n667), .B(n660), .ZN(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(G305), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n663), .B(n662), .ZN(n890) );
  XNOR2_X1 U747 ( .A(n664), .B(n890), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n665), .A2(G868), .ZN(n669) );
  INV_X1 U749 ( .A(G868), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(KEYINPUT85), .B(n670), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G69), .A2(G120), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT87), .B(n675), .Z(n676) );
  NOR2_X1 U761 ( .A1(G238), .A2(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G57), .A2(n677), .ZN(n825) );
  NAND2_X1 U763 ( .A1(n825), .A2(G567), .ZN(n683) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U766 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G96), .A2(n680), .ZN(n824) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n824), .ZN(n681) );
  XNOR2_X1 U769 ( .A(KEYINPUT86), .B(n681), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n826) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n826), .A2(n684), .ZN(n821) );
  NAND2_X1 U773 ( .A1(n821), .A2(G36), .ZN(G176) );
  XNOR2_X1 U774 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n771) );
  INV_X1 U776 ( .A(n771), .ZN(n685) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X1 U778 ( .A1(G1996), .A2(n714), .ZN(n687) );
  XNOR2_X1 U779 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n686) );
  XNOR2_X1 U780 ( .A(n687), .B(n686), .ZN(n691) );
  XOR2_X1 U781 ( .A(KEYINPUT98), .B(n688), .Z(n689) );
  NOR2_X1 U782 ( .A1(n932), .A2(n689), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n697) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT99), .ZN(n696) );
  NOR2_X1 U785 ( .A1(n714), .A2(G1348), .ZN(n694) );
  NOR2_X1 U786 ( .A1(G2067), .A2(n730), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n697), .A2(n912), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n714), .ZN(n702) );
  XOR2_X1 U792 ( .A(G1956), .B(KEYINPUT96), .Z(n990) );
  NOR2_X1 U793 ( .A1(n714), .A2(n990), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n712) );
  NOR2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U798 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n709) );
  XNOR2_X1 U799 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(KEYINPUT29), .B(n713), .ZN(n719) );
  NAND2_X1 U802 ( .A1(G1961), .A2(n730), .ZN(n716) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NAND2_X1 U804 ( .A1(n714), .A2(n944), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U806 ( .A1(G301), .A2(n720), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n717), .B(KEYINPUT94), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n729) );
  AND2_X1 U809 ( .A1(G301), .A2(n720), .ZN(n725) );
  NAND2_X1 U810 ( .A1(G8), .A2(n730), .ZN(n764) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n764), .ZN(n741) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n730), .ZN(n742) );
  NOR2_X1 U813 ( .A1(n741), .A2(n742), .ZN(n721) );
  NAND2_X1 U814 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n722), .ZN(n723) );
  NOR2_X1 U816 ( .A1(G168), .A2(n723), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT31), .B(n726), .ZN(n727) );
  XNOR2_X1 U819 ( .A(KEYINPUT100), .B(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n740) );
  OR2_X1 U821 ( .A1(n740), .A2(n514), .ZN(n738) );
  INV_X1 U822 ( .A(G8), .ZN(n736) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n764), .ZN(n732) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(KEYINPUT102), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n734), .A2(G303), .ZN(n735) );
  OR2_X1 U828 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U830 ( .A1(G8), .A2(n742), .ZN(n743) );
  AND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U832 ( .A(KEYINPUT101), .B(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n758) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n752), .A2(n748), .ZN(n925) );
  NAND2_X1 U837 ( .A1(n758), .A2(n925), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n917) );
  AND2_X1 U839 ( .A1(n750), .A2(n516), .ZN(n751) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n751), .ZN(n755) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n927) );
  NAND2_X1 U842 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n759), .A2(n764), .ZN(n766) );
  XNOR2_X1 U848 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(KEYINPUT92), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n762), .B(n761), .ZN(n763) );
  OR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U855 ( .A(n770), .B(n769), .ZN(n803) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n814) );
  NAND2_X1 U857 ( .A1(G116), .A2(n868), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G128), .A2(n869), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U860 ( .A(n775), .B(KEYINPUT35), .ZN(n780) );
  NAND2_X1 U861 ( .A1(n605), .A2(G104), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G140), .A2(n865), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U864 ( .A(KEYINPUT34), .B(n778), .Z(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U866 ( .A(n781), .B(KEYINPUT36), .Z(n880) );
  XNOR2_X1 U867 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  NOR2_X1 U868 ( .A1(n880), .A2(n811), .ZN(n971) );
  NAND2_X1 U869 ( .A1(n814), .A2(n971), .ZN(n809) );
  NAND2_X1 U870 ( .A1(G131), .A2(n865), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT90), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G95), .A2(n605), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U874 ( .A(KEYINPUT91), .B(n785), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n869), .A2(G119), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G107), .A2(n868), .ZN(n786) );
  AND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n883) );
  AND2_X1 U879 ( .A1(n883), .A2(G1991), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G117), .A2(n868), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G141), .A2(n865), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n605), .A2(G105), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G129), .A2(n869), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n875) );
  AND2_X1 U888 ( .A1(n875), .A2(G1996), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n959) );
  INV_X1 U890 ( .A(n814), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n959), .A2(n799), .ZN(n806) );
  INV_X1 U892 ( .A(n806), .ZN(n800) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n923) );
  NAND2_X1 U894 ( .A1(n923), .A2(n814), .ZN(n801) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n875), .ZN(n966) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n883), .ZN(n970) );
  NOR2_X1 U898 ( .A1(n804), .A2(n970), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n966), .A2(n807), .ZN(n808) );
  XNOR2_X1 U901 ( .A(KEYINPUT39), .B(n808), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n813) );
  AND2_X1 U903 ( .A1(n880), .A2(n811), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT104), .B(n812), .Z(n960) );
  NAND2_X1 U905 ( .A1(n813), .A2(n960), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U911 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G1), .A2(G3), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n823), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U915 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  INV_X1 U918 ( .A(G69), .ZN(G235) );
  NOR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U920 ( .A(G325), .ZN(G261) );
  INV_X1 U921 ( .A(n826), .ZN(G319) );
  XOR2_X1 U922 ( .A(G2096), .B(KEYINPUT43), .Z(n828) );
  XNOR2_X1 U923 ( .A(G2067), .B(G2678), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U925 ( .A(n829), .B(KEYINPUT110), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2072), .B(G2090), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(G2100), .Z(n833) );
  XNOR2_X1 U929 ( .A(G2084), .B(G2078), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U932 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n837) );
  XNOR2_X1 U933 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U935 ( .A(n838), .B(KEYINPUT113), .Z(n840) );
  XNOR2_X1 U936 ( .A(G1961), .B(G1971), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n848) );
  XOR2_X1 U938 ( .A(G1976), .B(G1956), .Z(n842) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(G2474), .B(G1981), .Z(n844) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G112), .A2(n868), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G100), .A2(n605), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n851), .B(KEYINPUT115), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G136), .A2(n865), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n869), .A2(G124), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n854), .Z(n855) );
  NOR2_X1 U954 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U955 ( .A1(G118), .A2(n868), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G130), .A2(n869), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U958 ( .A1(n605), .A2(G106), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G142), .A2(n865), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT116), .B(n862), .ZN(n863) );
  NOR2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n879) );
  XOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n877) );
  NAND2_X1 U965 ( .A1(n605), .A2(G103), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G115), .A2(n868), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G127), .A2(n869), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n961) );
  XOR2_X1 U973 ( .A(n875), .B(n961), .Z(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n882) );
  XOR2_X1 U976 ( .A(n880), .B(G162), .Z(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(n884) );
  XNOR2_X1 U978 ( .A(n884), .B(n883), .ZN(n886) );
  XNOR2_X1 U979 ( .A(G164), .B(G160), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n887), .B(n975), .ZN(n888) );
  NOR2_X1 U982 ( .A1(G37), .A2(n888), .ZN(n889) );
  XOR2_X1 U983 ( .A(KEYINPUT117), .B(n889), .Z(G395) );
  XNOR2_X1 U984 ( .A(G286), .B(n912), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n892), .B(G301), .ZN(n893) );
  NOR2_X1 U987 ( .A1(G37), .A2(n893), .ZN(G397) );
  XOR2_X1 U988 ( .A(G2438), .B(KEYINPUT106), .Z(n895) );
  XNOR2_X1 U989 ( .A(G2454), .B(G2435), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U991 ( .A(n896), .B(G2430), .Z(n898) );
  XNOR2_X1 U992 ( .A(G1341), .B(G1348), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U994 ( .A(G2446), .B(KEYINPUT107), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2451), .B(G2427), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U998 ( .A(KEYINPUT105), .B(G2443), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(n905), .A2(G14), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G301), .ZN(G171) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  INV_X1 U1010 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(G301), .B(G1961), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n912), .B(G1348), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT122), .B(n915), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(G1956), .B(G299), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT123), .B(n926), .ZN(n931) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n929), .B(KEYINPUT57), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G1341), .B(n932), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1029 ( .A(KEYINPUT56), .B(G16), .Z(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(KEYINPUT124), .B(n937), .Z(n989) );
  XNOR2_X1 U1032 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n982) );
  XOR2_X1 U1033 ( .A(G25), .B(G1991), .Z(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(n941), .B(KEYINPUT121), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G1996), .B(G32), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G27), .B(n944), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n949), .B(KEYINPUT53), .ZN(n952) );
  XOR2_X1 U1045 ( .A(G2084), .B(G34), .Z(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n950), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(n982), .B(n955), .Z(n957) );
  INV_X1 U1051 ( .A(G29), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G11), .ZN(n987) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n980) );
  XOR2_X1 U1055 ( .A(G2072), .B(n961), .Z(n963) );
  XOR2_X1 U1056 ( .A(G164), .B(G2078), .Z(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT50), .B(n964), .Z(n969) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT51), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n978) );
  XNOR2_X1 U1063 ( .A(G160), .B(G2084), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n976), .B(KEYINPUT118), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(KEYINPUT52), .B(n981), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n984), .A2(G29), .ZN(n985) );
  XOR2_X1 U1073 ( .A(KEYINPUT120), .B(n985), .Z(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n1016) );
  XNOR2_X1 U1076 ( .A(n990), .B(G20), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(G1341), .B(G19), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G6), .B(G1981), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1081 ( .A(KEYINPUT59), .B(G1348), .Z(n995) );
  XNOR2_X1 U1082 ( .A(G4), .B(n995), .ZN(n996) );
  NOR2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT60), .B(n998), .ZN(n1011) );
  XOR2_X1 U1085 ( .A(G1961), .B(G5), .Z(n1006) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1976), .B(G23), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(n1001), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(G21), .B(G1966), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT125), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(KEYINPUT61), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1013), .Z(n1014) );
  NOR2_X1 U1100 ( .A1(G16), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1017), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

