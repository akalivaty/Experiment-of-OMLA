//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT76), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n187), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n188), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n196), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n199));
  OAI211_X1 g013(.A(G119), .B(new_n187), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT75), .B1(new_n201), .B2(G110), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n203));
  INV_X1    g017(.A(G110), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n197), .A2(new_n200), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n194), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(KEYINPUT78), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n208), .A2(new_n210), .A3(new_n216), .A4(KEYINPUT16), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT16), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT74), .B1(new_n208), .B2(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT77), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(KEYINPUT74), .C1(KEYINPUT16), .C2(new_n208), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n212), .B1(new_n224), .B2(new_n217), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n206), .A2(new_n215), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n201), .A2(G110), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n212), .A3(new_n217), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI221_X1 g045(.A(new_n229), .B1(new_n191), .B2(new_n192), .C1(new_n231), .C2(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n232), .A3(KEYINPUT80), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT79), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G137), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT80), .B1(new_n228), .B2(new_n232), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI211_X1 g056(.A(KEYINPUT80), .B(new_n239), .C1(new_n228), .C2(new_n232), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G217), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(G234), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G902), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  AOI21_X1  g066(.A(G902), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n241), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n233), .A3(new_n239), .ZN(new_n256));
  INV_X1    g070(.A(new_n243), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n251), .A2(new_n252), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n248), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(new_n242), .B2(new_n243), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n250), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n212), .A2(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G137), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT11), .A3(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(G137), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G131), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n284), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(new_n278), .A3(new_n280), .A4(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n275), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n283), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n283), .B1(G134), .B2(new_n279), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n273), .A2(new_n294), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n269), .A2(new_n187), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n212), .A2(G143), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n289), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT30), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n290), .A2(new_n307), .A3(new_n292), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(new_n302), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT67), .B1(new_n275), .B2(new_n288), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n305), .B1(new_n312), .B2(KEYINPUT30), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G113), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G116), .B(G119), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n189), .A2(G116), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G113), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT66), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n265), .B1(new_n313), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n289), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n275), .A2(new_n288), .A3(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n309), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT69), .B(new_n331), .C1(new_n337), .C2(new_n305), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n309), .B(new_n329), .C1(new_n310), .C2(new_n311), .ZN(new_n339));
  INV_X1    g153(.A(G237), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n234), .A3(G210), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n341), .B(KEYINPUT27), .Z(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G101), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND4_X1  g158(.A1(new_n330), .A2(new_n338), .A3(new_n339), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT31), .ZN(new_n346));
  INV_X1    g160(.A(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n312), .A2(KEYINPUT30), .ZN(new_n348));
  INV_X1    g162(.A(new_n305), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n329), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n350), .B2(KEYINPUT69), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n344), .A4(new_n330), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n309), .A2(new_n329), .A3(new_n289), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n355), .B1(new_n354), .B2(new_n356), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n304), .A2(new_n331), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n304), .A2(KEYINPUT70), .A3(new_n331), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n339), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n344), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n346), .A2(new_n353), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT72), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n375), .B(KEYINPUT32), .C1(new_n370), .C2(new_n371), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n366), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n354), .A2(new_n356), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n357), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n312), .A2(new_n331), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n356), .B1(new_n384), .B2(new_n339), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT29), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n386), .A3(new_n344), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n351), .A2(new_n379), .A3(new_n368), .A4(new_n330), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n247), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G472), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n264), .B1(new_n377), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(KEYINPUT3), .A2(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(KEYINPUT3), .A2(G107), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(G104), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(KEYINPUT83), .A2(G104), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT83), .A2(G104), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(G104), .B2(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n295), .B(new_n296), .C1(new_n298), .C2(new_n267), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n410), .A2(new_n411), .B1(new_n412), .B2(new_n302), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n272), .A2(new_n274), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  INV_X1    g229(.A(new_n400), .ZN(new_n416));
  NOR2_X1   g230(.A1(KEYINPUT83), .A2(G104), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n416), .A2(new_n394), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n397), .A2(new_n398), .A3(G104), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT3), .A2(G107), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n415), .B(G101), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n395), .A2(new_n401), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n425), .A2(KEYINPUT85), .A3(new_n415), .A4(G101), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n414), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G101), .B1(new_n418), .B2(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT84), .B(G101), .C1(new_n418), .C2(new_n421), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n430), .A2(KEYINPUT4), .A3(new_n431), .A4(new_n403), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n288), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n413), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n408), .A2(KEYINPUT86), .A3(new_n302), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n434), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n410), .B(KEYINPUT86), .C1(new_n302), .C2(new_n408), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT12), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT12), .B1(new_n437), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G140), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT82), .ZN(new_n443));
  INV_X1    g257(.A(G227), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G953), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n443), .B(new_n445), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n413), .A2(new_n433), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n413), .A2(new_n433), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n288), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n435), .A2(new_n446), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n441), .A2(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G469), .B1(new_n454), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n446), .B1(new_n452), .B2(new_n435), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n439), .A2(new_n440), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n435), .A2(new_n446), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n456), .B(new_n247), .C1(new_n457), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT9), .B(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT92), .B(G143), .ZN(new_n467));
  INV_X1    g281(.A(G214), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n468), .A2(G237), .A3(G953), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n266), .A2(KEYINPUT92), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n283), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n473), .A2(KEYINPUT93), .A3(new_n283), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n469), .B1(new_n477), .B2(G143), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n469), .B2(new_n467), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n479), .B2(G131), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n466), .B(new_n474), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n222), .A2(new_n230), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(G131), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n476), .A3(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(KEYINPUT17), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT94), .B1(new_n231), .B2(new_n225), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n481), .A2(new_n483), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(G104), .Z(new_n491));
  INV_X1    g305(.A(KEYINPUT18), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n473), .B1(new_n492), .B2(new_n283), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n211), .A2(new_n212), .ZN(new_n494));
  OAI221_X1 g308(.A(new_n493), .B1(new_n492), .B2(new_n484), .C1(new_n214), .C2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n489), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n491), .B1(new_n489), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n247), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT96), .B(G475), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n211), .B(KEYINPUT19), .Z(new_n502));
  OAI211_X1 g316(.A(new_n223), .B(new_n227), .C1(G146), .C2(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n485), .A2(new_n486), .B1(new_n283), .B2(new_n473), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n495), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n491), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n489), .A2(new_n491), .A3(new_n495), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT95), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n501), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI211_X1 g327(.A(KEYINPUT20), .B(new_n511), .C1(new_n507), .C2(new_n508), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n500), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(G234), .A2(G237), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n517), .A2(G952), .A3(new_n234), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n517), .A2(G902), .A3(G953), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT21), .B(G898), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n323), .A2(G122), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT99), .B1(new_n523), .B2(KEYINPUT14), .ZN(new_n524));
  INV_X1    g338(.A(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G116), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(KEYINPUT14), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n523), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g343(.A(G107), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT97), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT97), .B1(new_n523), .B2(new_n526), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n398), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G128), .B(G143), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n277), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n277), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n266), .A2(KEYINPUT13), .A3(G128), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT98), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n187), .B2(G143), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n544), .C1(G128), .C2(new_n266), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n541), .A2(KEYINPUT98), .ZN(new_n546));
  OAI21_X1  g360(.A(G134), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n534), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n532), .A2(new_n398), .A3(new_n533), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n540), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n537), .A2(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n539), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n463), .A2(new_n246), .A3(G953), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n539), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n247), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n558), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n516), .A2(new_n522), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT88), .B1(new_n322), .B2(KEYINPUT5), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT5), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n189), .A4(G116), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n565), .A2(new_n566), .A3(G113), .A4(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n325), .A2(new_n326), .A3(new_n321), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT66), .B1(new_n318), .B2(new_n319), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n407), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n426), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n402), .B1(new_n395), .B2(new_n401), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT85), .B1(new_n577), .B2(new_n415), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n331), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(KEYINPUT84), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n575), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT89), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G122), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n329), .B1(new_n424), .B2(new_n426), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n574), .B1(new_n588), .B2(new_n432), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT89), .B1(new_n589), .B2(new_n585), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT6), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n589), .B2(new_n585), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n302), .A2(G125), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n414), .A2(G125), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G224), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n589), .A2(new_n585), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  NOR4_X1   g416(.A1(new_n589), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n585), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n593), .B(new_n599), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n596), .A2(new_n605), .A3(new_n598), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n585), .B(KEYINPUT8), .Z(new_n607));
  NAND2_X1  g421(.A1(new_n573), .A2(new_n407), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n575), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n598), .A2(new_n605), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n594), .B2(new_n595), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n589), .A2(new_n585), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(G210), .B1(G237), .B2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n604), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n604), .B2(new_n614), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G214), .B1(G237), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n564), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n604), .A2(new_n614), .ZN(new_n623));
  INV_X1    g437(.A(new_n615), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n616), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(KEYINPUT91), .A3(new_n620), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n465), .B(new_n563), .C1(new_n622), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n392), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  NOR2_X1   g444(.A1(new_n465), .A2(new_n264), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n370), .A2(new_n247), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n370), .B2(new_n247), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n631), .A2(new_n634), .A3(new_n372), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n639));
  INV_X1    g453(.A(new_n637), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n372), .B1(new_n635), .B2(new_n636), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n631), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT104), .B1(new_n623), .B2(new_n624), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n647), .B(new_n615), .C1(new_n604), .C2(new_n614), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n616), .A2(KEYINPUT103), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n604), .A2(new_n651), .A3(new_n614), .A4(new_n615), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n621), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n555), .A2(new_n655), .A3(new_n556), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n555), .B2(new_n556), .ZN(new_n657));
  OAI211_X1 g471(.A(G478), .B(new_n247), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT105), .B(G478), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n558), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n516), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n654), .A2(new_n522), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n645), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT34), .B(G104), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  XNOR2_X1  g481(.A(new_n521), .B(KEYINPUT106), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n515), .A2(new_n562), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n654), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n228), .A2(new_n232), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n239), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n249), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n261), .B2(new_n263), .ZN(new_n678));
  INV_X1    g492(.A(new_n464), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n455), .B2(new_n461), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n563), .B(new_n681), .C1(new_n622), .C2(new_n627), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n642), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT37), .B(G110), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT107), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n683), .B(new_n685), .ZN(G12));
  AOI21_X1  g500(.A(new_n681), .B1(new_n377), .B2(new_n391), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n519), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n518), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n515), .A2(new_n562), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n654), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n625), .A2(new_n647), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n618), .A2(KEYINPUT104), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n653), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(KEYINPUT108), .A2(new_n695), .A3(new_n620), .A4(new_n691), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n687), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT109), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n620), .A3(new_n691), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n654), .A2(KEYINPUT108), .A3(new_n691), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n687), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  NAND2_X1  g521(.A1(new_n372), .A2(new_n373), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n375), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n368), .B1(new_n351), .B2(new_n330), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n384), .A2(new_n339), .A3(new_n368), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n247), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n378), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT32), .B1(new_n370), .B2(new_n371), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT72), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n709), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n678), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n690), .B(KEYINPUT39), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n680), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT40), .Z(new_n722));
  NOR3_X1   g536(.A1(new_n516), .A2(new_n621), .A3(new_n562), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT38), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n626), .B(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n719), .A2(new_n722), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G143), .ZN(G45));
  NAND3_X1  g542(.A1(new_n709), .A2(new_n391), .A3(new_n716), .ZN(new_n729));
  INV_X1    g543(.A(new_n690), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n515), .A2(new_n661), .A3(new_n730), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n621), .B(new_n731), .C1(new_n649), .C2(new_n653), .ZN(new_n732));
  INV_X1    g546(.A(new_n681), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  OAI21_X1  g549(.A(new_n247), .B1(new_n457), .B2(new_n460), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n461), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n679), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n392), .A2(new_n664), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND3_X1  g556(.A1(new_n392), .A2(new_n670), .A3(new_n739), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  INV_X1    g558(.A(new_n248), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n262), .B2(new_n259), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n258), .A2(new_n260), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n746), .A2(new_n747), .B1(new_n249), .B2(new_n676), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n563), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n654), .A2(new_n739), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n729), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  AND4_X1   g566(.A1(new_n695), .A2(new_n739), .A3(new_n668), .A4(new_n723), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n368), .B1(new_n383), .B2(new_n385), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n346), .A2(new_n353), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n371), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n635), .A3(new_n264), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT110), .B(G122), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G24));
  NOR3_X1   g574(.A1(new_n756), .A2(new_n748), .A3(new_n635), .ZN(new_n761));
  INV_X1    g575(.A(new_n731), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n654), .A3(new_n762), .A4(new_n739), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  INV_X1    g578(.A(new_n264), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n619), .A2(new_n620), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n465), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n729), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n378), .A2(new_n390), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n765), .B1(new_n770), .B2(new_n715), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n626), .A2(new_n621), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n762), .A3(new_n680), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND4_X1  g590(.A1(new_n729), .A2(new_n765), .A3(new_n691), .A4(new_n767), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n781));
  OAI22_X1  g595(.A1(new_n662), .A2(new_n515), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n516), .A2(new_n661), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(new_n781), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n678), .C1(new_n640), .C2(new_n641), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n772), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n786), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n454), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n454), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n461), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n464), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n720), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NOR4_X1   g618(.A1(new_n729), .A2(new_n765), .A3(new_n731), .A4(new_n766), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT114), .Z(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(KEYINPUT113), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n806), .B(new_n810), .C1(new_n801), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n516), .A2(new_n562), .A3(new_n730), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n766), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n687), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n729), .A2(new_n816), .A3(new_n733), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n622), .A2(new_n627), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n663), .A2(new_n669), .ZN(new_n822));
  INV_X1    g636(.A(new_n668), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n639), .A2(new_n644), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n761), .A2(new_n767), .A3(new_n762), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n777), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n642), .A2(new_n682), .B1(new_n392), .B2(new_n628), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n750), .A2(new_n729), .B1(new_n753), .B2(new_n757), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n775), .A2(new_n830), .A3(new_n740), .A4(new_n743), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n695), .A2(new_n723), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n465), .A2(new_n690), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n717), .A2(new_n833), .A3(new_n748), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(new_n734), .A3(new_n763), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n706), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n734), .A3(new_n763), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n838), .B(new_n839), .C1(new_n698), .C2(new_n705), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n832), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n703), .A2(new_n704), .A3(new_n687), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n704), .B1(new_n703), .B2(new_n687), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n838), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  OAI211_X1 g661(.A(KEYINPUT52), .B(new_n836), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n837), .A2(KEYINPUT116), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n852), .A3(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n855), .B(new_n831), .C1(KEYINPUT118), .C2(new_n829), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n849), .A3(new_n850), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n841), .A2(new_n855), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n842), .A2(new_n852), .A3(new_n862), .A4(KEYINPUT54), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n757), .A2(new_n784), .A3(new_n518), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n725), .A2(new_n621), .A3(new_n739), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n739), .A2(new_n518), .A3(new_n772), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n761), .A3(new_n784), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n718), .A2(new_n765), .A3(new_n870), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n516), .A3(new_n662), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n869), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT120), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n737), .A2(new_n679), .A3(new_n461), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n801), .A2(new_n809), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n801), .A2(new_n811), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n864), .A2(new_n766), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n869), .A2(new_n873), .A3(new_n882), .A4(new_n871), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(KEYINPUT51), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n771), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n870), .A2(new_n885), .A3(new_n784), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT48), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n872), .A2(new_n663), .ZN(new_n888));
  INV_X1    g702(.A(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n864), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n654), .A2(new_n739), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n889), .B(G953), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n887), .A2(new_n895), .A3(new_n888), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT119), .B1(new_n877), .B2(new_n878), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n810), .B(new_n899), .C1(new_n801), .C2(new_n811), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n876), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n874), .B1(new_n901), .B2(new_n880), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n884), .B(new_n897), .C1(new_n902), .C2(KEYINPUT51), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n854), .A2(new_n861), .A3(new_n863), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n889), .A2(new_n234), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n783), .A2(new_n679), .A3(new_n621), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n765), .C1(KEYINPUT49), .C2(new_n738), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(KEYINPUT49), .B2(new_n738), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n718), .A3(new_n725), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n234), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n247), .B1(new_n858), .B2(new_n860), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n593), .B1(new_n602), .B2(new_n603), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n599), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n920), .B2(new_n923), .ZN(G51));
  NAND2_X1  g739(.A1(new_n858), .A2(new_n860), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n861), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n795), .B(KEYINPUT57), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n457), .B2(new_n460), .ZN(new_n931));
  INV_X1    g745(.A(new_n794), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n917), .B1(new_n931), .B2(new_n933), .ZN(G54));
  AND2_X1   g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n919), .A2(new_n509), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n509), .B1(new_n919), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n917), .ZN(G60));
  OR2_X1    g752(.A1(new_n656), .A2(new_n657), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n928), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n854), .A2(new_n861), .A3(new_n863), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n944), .B2(new_n942), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n945), .A3(new_n917), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n858), .B2(new_n860), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n676), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n918), .C1(new_n245), .C2(new_n951), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT61), .B1(new_n952), .B2(KEYINPUT125), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  OAI21_X1  g769(.A(G953), .B1(new_n520), .B2(new_n597), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n830), .A2(new_n740), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n743), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n825), .A2(new_n828), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n960), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n921), .B1(G898), .B2(new_n234), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  AND3_X1   g777(.A1(new_n706), .A2(new_n734), .A3(new_n763), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n727), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT127), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n822), .A2(new_n721), .A3(new_n766), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n392), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n812), .A2(new_n803), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(KEYINPUT62), .B2(new_n965), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n502), .B(KEYINPUT126), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n313), .B(new_n973), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n802), .A2(new_n833), .A3(new_n885), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n775), .A2(new_n812), .A3(new_n777), .A4(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n803), .A3(new_n964), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(G953), .B1(new_n980), .B2(new_n974), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n974), .A2(G227), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n688), .B(new_n234), .C1(new_n975), .C2(new_n444), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n976), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n960), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n351), .A2(new_n368), .A3(new_n330), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n986), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n989), .A2(new_n710), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n842), .A2(new_n852), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n918), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n972), .B2(new_n987), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n710), .ZN(G57));
endmodule


