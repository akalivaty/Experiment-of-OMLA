//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n188), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT75), .B(KEYINPUT27), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n192), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n195), .A2(KEYINPUT67), .A3(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  OR3_X1    g011(.A1(new_n197), .A2(KEYINPUT68), .A3(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT67), .B1(new_n195), .B2(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n197), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n197), .A3(G134), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT69), .B(KEYINPUT1), .C1(new_n213), .C2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G128), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(G143), .B(G146), .Z(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n219), .A2(KEYINPUT1), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT73), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n214), .B2(new_n215), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n217), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n219), .A2(KEYINPUT1), .A3(new_n221), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT73), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n212), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT2), .A2(G113), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT71), .B1(KEYINPUT2), .B2(G113), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(KEYINPUT2), .B2(G113), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(new_n235), .B2(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT65), .B1(new_n208), .B2(new_n209), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n206), .B1(G134), .B2(new_n197), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n195), .A2(KEYINPUT11), .A3(G137), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n200), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(KEYINPUT65), .A3(G131), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n219), .A2(KEYINPUT64), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n224), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n230), .A2(new_n242), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(KEYINPUT78), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n242), .B1(new_n230), .B2(new_n256), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n230), .A2(KEYINPUT74), .A3(new_n242), .A4(new_n256), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n259), .B(new_n262), .C1(new_n267), .C2(new_n258), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n194), .B1(new_n268), .B2(KEYINPUT29), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n256), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n220), .A2(new_n222), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n212), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n248), .A2(KEYINPUT66), .A3(new_n249), .A4(new_n255), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n265), .A2(new_n266), .B1(new_n241), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT77), .B(KEYINPUT28), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n270), .B(new_n260), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n230), .A2(new_n256), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n276), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n283), .A2(new_n241), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(new_n266), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n287), .A2(new_n194), .A3(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n269), .A2(new_n279), .B1(new_n270), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT79), .B(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n187), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n260), .B1(new_n277), .B2(new_n278), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n194), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n194), .B1(new_n265), .B2(new_n266), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n287), .B2(new_n297), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n287), .A2(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n300), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n295), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n293), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n310));
  INV_X1    g124(.A(new_n306), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n302), .A2(KEYINPUT76), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT31), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n303), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(new_n295), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n316), .B2(KEYINPUT32), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n314), .A2(new_n303), .B1(new_n194), .B2(new_n294), .ZN(new_n318));
  NOR4_X1   g132(.A1(new_n318), .A2(KEYINPUT80), .A3(new_n308), .A4(new_n311), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n309), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n292), .B2(G234), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G128), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT23), .B1(new_n221), .B2(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n324), .B(new_n331), .C1(new_n327), .C2(KEYINPUT82), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G110), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n221), .A2(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT24), .B(G110), .Z(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT83), .ZN(new_n341));
  INV_X1    g155(.A(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(KEYINPUT16), .B2(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n347), .A2(new_n342), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(G146), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n337), .B2(new_n338), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n334), .B2(new_n333), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n353), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n292), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT25), .B1(new_n357), .B2(new_n292), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n322), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n322), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n320), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT80), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n316), .A2(new_n310), .A3(KEYINPUT32), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n365), .B1(new_n373), .B2(new_n309), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT84), .ZN(new_n375));
  INV_X1    g189(.A(G475), .ZN(new_n376));
  INV_X1    g190(.A(G902), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT96), .B(G104), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(G143), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT95), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n340), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n341), .B2(new_n386), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n342), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n348), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n383), .B(new_n391), .Z(new_n392));
  INV_X1    g206(.A(new_n343), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n340), .A2(new_n342), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT94), .Z(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n381), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n350), .A2(KEYINPUT98), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n347), .B(new_n342), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT98), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  OR3_X1    g216(.A1(new_n383), .A2(new_n402), .A3(new_n209), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n384), .A2(new_n402), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n398), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n380), .B(KEYINPUT97), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n405), .A2(new_n396), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n376), .B(new_n377), .C1(new_n397), .C2(new_n407), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(KEYINPUT20), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(KEYINPUT20), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n381), .B1(new_n405), .B2(new_n396), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n377), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n409), .A2(new_n410), .B1(G475), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n190), .A2(G952), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(G234), .B2(G237), .ZN(new_n415));
  NAND2_X1  g229(.A1(G234), .A2(G237), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n291), .A2(G953), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT21), .B(G898), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n415), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n221), .A2(G143), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT99), .Z(new_n425));
  NOR2_X1   g239(.A1(new_n213), .A2(G128), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n423), .B2(KEYINPUT13), .ZN(new_n428));
  OAI21_X1  g242(.A(G134), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n423), .A2(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n195), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G122), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n429), .B(new_n431), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n430), .B(new_n195), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT100), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT101), .ZN(new_n439));
  INV_X1    g253(.A(G116), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n440), .A2(KEYINPUT14), .A3(G122), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n432), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n434), .B1(new_n443), .B2(G107), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n438), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n439), .B1(new_n438), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n436), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT9), .B(G234), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT85), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G217), .A3(new_n190), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n450), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n436), .B(new_n452), .C1(new_n445), .C2(new_n446), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n292), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n455), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n413), .A2(new_n422), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT102), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n190), .A2(G227), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n345), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT87), .B(G110), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n214), .A2(G128), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n222), .B1(new_n467), .B2(new_n224), .ZN(new_n468));
  INV_X1    g282(.A(G101), .ZN(new_n469));
  INV_X1    g283(.A(G104), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n470), .A2(KEYINPUT3), .A3(G107), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G104), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n475), .B2(G107), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n474), .A3(new_n433), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT3), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n477), .B2(KEYINPUT3), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n469), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(G104), .B2(new_n433), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G101), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n468), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT10), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT10), .B1(new_n223), .B2(new_n229), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n483), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G101), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n481), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n494), .A3(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n255), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT90), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n493), .A2(new_n498), .A3(new_n255), .A4(new_n495), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n487), .B(new_n490), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n248), .A2(new_n249), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n466), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n499), .ZN(new_n503));
  INV_X1    g317(.A(new_n490), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n486), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n503), .A2(new_n501), .A3(new_n486), .A4(new_n504), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n226), .A2(new_n227), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n489), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT91), .A3(new_n484), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n489), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n511), .A2(KEYINPUT12), .A3(new_n506), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n502), .A2(new_n507), .B1(new_n519), .B2(new_n466), .ZN(new_n520));
  OAI21_X1  g334(.A(G469), .B1(new_n520), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(G469), .ZN(new_n522));
  INV_X1    g336(.A(new_n466), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n507), .B2(new_n508), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n508), .A2(new_n523), .A3(new_n518), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n522), .B(new_n292), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n449), .A2(new_n377), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G221), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT86), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(G110), .B(G122), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n493), .A2(new_n495), .A3(new_n241), .ZN(new_n534));
  INV_X1    g348(.A(G113), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n440), .A2(KEYINPUT5), .A3(G119), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n535), .B(new_n536), .C1(new_n237), .C2(KEYINPUT5), .ZN(new_n537));
  INV_X1    g351(.A(new_n240), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n238), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n481), .A3(new_n483), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n481), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n495), .A2(new_n241), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n540), .B(new_n533), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n534), .A2(KEYINPUT92), .A3(new_n540), .A4(new_n533), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G125), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n273), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n255), .A2(G125), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G224), .A3(new_n190), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n190), .A2(G224), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT7), .B1(new_n190), .B2(G224), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n559), .B(new_n562), .Z(new_n563));
  XOR2_X1   g377(.A(new_n539), .B(new_n489), .Z(new_n564));
  XOR2_X1   g378(.A(new_n532), .B(KEYINPUT8), .Z(new_n565));
  AOI22_X1  g379(.A1(new_n547), .A2(new_n548), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G210), .B1(G237), .B2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n569), .A3(new_n567), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT93), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(KEYINPUT93), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G214), .B1(G237), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR4_X1   g392(.A1(new_n462), .A2(new_n531), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n369), .A2(new_n375), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT103), .B(G101), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G3));
  OAI21_X1  g396(.A(G472), .B1(new_n318), .B2(new_n291), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n307), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n531), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n366), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n561), .A2(new_n569), .A3(new_n567), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n569), .B1(new_n561), .B2(new_n567), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n577), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT105), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n454), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n451), .A2(KEYINPUT33), .A3(new_n453), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(G478), .A3(new_n292), .A4(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n455), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n598), .B1(G478), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n412), .A2(G475), .ZN(new_n601));
  INV_X1    g415(.A(new_n410), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n408), .A2(KEYINPUT20), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n607), .B(new_n577), .C1(new_n591), .C2(new_n592), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n422), .A2(new_n594), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NOR2_X1   g427(.A1(new_n604), .A2(new_n459), .ZN(new_n614));
  AND4_X1   g428(.A1(new_n422), .A2(new_n594), .A3(new_n608), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n590), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT35), .B(G107), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n356), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n353), .B(new_n621), .Z(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n363), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n362), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n579), .A2(new_n588), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n530), .A3(new_n527), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n373), .B2(new_n309), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n594), .A2(new_n608), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n415), .B(KEYINPUT106), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n417), .A2(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n604), .A2(new_n459), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NOR2_X1   g452(.A1(new_n413), .A2(new_n459), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n634), .B(KEYINPUT39), .Z(new_n640));
  NOR2_X1   g454(.A1(new_n531), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n639), .B1(new_n642), .B2(KEYINPUT40), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n307), .A2(new_n308), .ZN(new_n644));
  INV_X1    g458(.A(new_n194), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n267), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n312), .B2(new_n313), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n647), .B2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n373), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT107), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n373), .A2(new_n651), .A3(new_n644), .A4(new_n648), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n643), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n624), .A2(new_n578), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n576), .B(KEYINPUT38), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  NOR2_X1   g473(.A1(new_n605), .A2(new_n635), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n629), .A2(new_n630), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  OAI21_X1  g476(.A(new_n292), .B1(new_n524), .B2(new_n525), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G469), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n529), .A3(new_n526), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n609), .A2(new_n320), .A3(new_n366), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n615), .A2(new_n320), .A3(new_n366), .A4(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  NAND4_X1  g484(.A1(new_n594), .A2(new_n665), .A3(new_n608), .A4(new_n624), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n462), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n320), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G119), .ZN(G21));
  AND3_X1   g489(.A1(new_n594), .A2(new_n608), .A3(new_n639), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n268), .A2(new_n194), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n315), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n306), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n314), .A2(new_n303), .B1(new_n194), .B2(new_n268), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT108), .B1(new_n681), .B2(new_n311), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n366), .A2(new_n680), .A3(new_n583), .A4(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n676), .A2(new_n683), .A3(new_n422), .A4(new_n665), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  AND3_X1   g499(.A1(new_n680), .A2(new_n583), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n672), .A2(new_n660), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G125), .ZN(G27));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n689));
  INV_X1    g503(.A(new_n529), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n521), .B2(new_n526), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT93), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n591), .B2(new_n592), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n693), .A3(new_n577), .A4(new_n574), .ZN(new_n694));
  INV_X1    g508(.A(new_n660), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT42), .B1(new_n374), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n309), .A2(new_n370), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n366), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n689), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n576), .A2(new_n577), .A3(new_n660), .A4(new_n691), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n367), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(KEYINPUT109), .B(new_n699), .C1(new_n703), .C2(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  INV_X1    g520(.A(new_n694), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n320), .A2(new_n366), .A3(new_n636), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  NOR3_X1   g523(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n413), .B2(KEYINPUT110), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n413), .A2(new_n600), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n413), .B(new_n600), .C1(KEYINPUT110), .C2(KEYINPUT43), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n587), .A2(new_n624), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n520), .A2(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n520), .A2(KEYINPUT45), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(G469), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(G469), .A2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n526), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT46), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n529), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(new_n640), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n716), .A2(new_n717), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT111), .B(new_n710), .C1(new_n716), .C2(new_n717), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n720), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  XNOR2_X1  g548(.A(new_n728), .B(KEYINPUT47), .ZN(new_n735));
  INV_X1    g549(.A(new_n710), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n366), .A3(new_n695), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n735), .A2(new_n320), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n345), .ZN(G42));
  INV_X1    g554(.A(new_n715), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n366), .A2(new_n680), .A3(new_n583), .A4(new_n682), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n632), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n630), .A3(new_n665), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n710), .A2(new_n665), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n366), .A2(new_n415), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n650), .A2(new_n745), .A3(new_n652), .A4(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n604), .A3(new_n600), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n664), .A2(new_n526), .ZN(new_n749));
  INV_X1    g563(.A(new_n530), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n736), .B1(new_n735), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n752), .B2(new_n743), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n743), .A2(new_n656), .A3(new_n578), .A4(new_n665), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT117), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n743), .A2(new_n656), .A3(new_n578), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT50), .A4(new_n665), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n754), .A2(new_n760), .A3(new_n755), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n754), .B2(new_n755), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n756), .B(new_n759), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n583), .A2(new_n680), .A3(new_n682), .A4(new_n624), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n745), .A2(new_n631), .A3(new_n715), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n753), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n414), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n747), .A2(new_n605), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n753), .A2(new_n763), .A3(KEYINPUT51), .A4(new_n765), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n744), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n455), .B(new_n457), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n604), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n693), .A2(new_n577), .A3(new_n574), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n635), .ZN(new_n775));
  INV_X1    g589(.A(new_n628), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n320), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n696), .A2(new_n764), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n708), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT113), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n708), .A2(new_n777), .A3(new_n781), .A4(new_n778), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n701), .A2(new_n704), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n606), .A2(new_n614), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n784), .A2(new_n576), .A3(new_n578), .A4(new_n421), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n588), .A2(new_n785), .A3(new_n589), .A4(new_n366), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n580), .A2(new_n625), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n666), .A2(new_n669), .A3(new_n674), .A4(new_n684), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n671), .A2(new_n462), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n594), .A2(new_n665), .A3(new_n608), .A4(new_n639), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n421), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n320), .A2(new_n792), .B1(new_n794), .B2(new_n683), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT112), .A3(new_n666), .A4(new_n669), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n783), .A2(new_n788), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n362), .A2(new_n623), .A3(new_n634), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n676), .A2(new_n691), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n800), .B(new_n801), .C1(new_n650), .C2(new_n652), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n637), .A2(new_n661), .A3(new_n687), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT114), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n799), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n802), .B2(new_n803), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n650), .A2(new_n652), .ZN(new_n810));
  INV_X1    g624(.A(new_n800), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n676), .A3(new_n691), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n637), .A2(new_n661), .A3(new_n687), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n805), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n798), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n808), .A2(KEYINPUT54), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n798), .B2(new_n815), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n666), .A2(new_n669), .A3(new_n674), .A4(new_n684), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n629), .A2(new_n775), .B1(new_n696), .B2(new_n764), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n781), .B1(new_n822), .B2(new_n708), .ZN(new_n823));
  INV_X1    g637(.A(new_n782), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n580), .A2(new_n625), .A3(new_n786), .A4(KEYINPUT53), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n699), .B1(new_n703), .B2(KEYINPUT42), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n806), .A3(new_n807), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n819), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n819), .A2(new_n820), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n771), .A2(new_n817), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n745), .A2(new_n631), .A3(new_n715), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n698), .A2(new_n366), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT48), .B1(new_n839), .B2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n840), .B(new_n841), .Z(new_n842));
  OAI22_X1  g656(.A1(new_n835), .A2(new_n842), .B1(G952), .B2(G953), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n750), .B1(new_n749), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n656), .A2(new_n577), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n366), .B1(new_n749), .B2(new_n844), .ZN(new_n847));
  OR4_X1    g661(.A1(new_n810), .A2(new_n846), .A3(new_n712), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(G75));
  XNOR2_X1  g663(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n292), .B(new_n569), .C1(new_n819), .C2(new_n829), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n551), .B(new_n559), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(KEYINPUT56), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n819), .A2(new_n829), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n291), .A3(new_n570), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n850), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n190), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n852), .B1(new_n851), .B2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n857), .A3(new_n854), .ZN(new_n863));
  INV_X1    g677(.A(new_n850), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n859), .A2(new_n861), .A3(new_n865), .ZN(G51));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n292), .B(new_n723), .C1(new_n819), .C2(new_n829), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n724), .B(KEYINPUT57), .Z(new_n869));
  AOI21_X1  g683(.A(new_n820), .B1(new_n819), .B2(new_n829), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n830), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n524), .ZN(new_n872));
  INV_X1    g686(.A(new_n525), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n868), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n867), .B1(new_n875), .B2(new_n860), .ZN(new_n876));
  INV_X1    g690(.A(new_n874), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n833), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n879), .B2(new_n869), .ZN(new_n880));
  OAI211_X1 g694(.A(KEYINPUT120), .B(new_n861), .C1(new_n880), .C2(new_n868), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n881), .ZN(G54));
  OR2_X1    g696(.A1(new_n397), .A2(new_n407), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n855), .A2(new_n291), .ZN(new_n885));
  AND3_X1   g699(.A1(KEYINPUT121), .A2(KEYINPUT58), .A3(G475), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(KEYINPUT58), .B2(G475), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR4_X1    g703(.A1(new_n884), .A2(new_n885), .A3(new_n888), .A4(new_n886), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n861), .ZN(G60));
  AND2_X1   g705(.A1(new_n596), .A2(new_n597), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n832), .A2(new_n834), .A3(new_n817), .ZN(new_n893));
  NAND2_X1  g707(.A1(G478), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT59), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n879), .A2(new_n892), .A3(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n898), .A3(new_n860), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n855), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n357), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n855), .A2(new_n622), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n861), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT61), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT61), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(G66));
  INV_X1    g724(.A(G224), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n420), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n787), .B1(new_n791), .B2(new_n796), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(G953), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  OAI221_X1 g729(.A(new_n542), .B1(G898), .B2(new_n190), .C1(new_n549), .C2(new_n550), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(G69));
  NAND3_X1  g731(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(new_n388), .Z(new_n919));
  NAND2_X1  g733(.A1(G900), .A2(G953), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n720), .A2(new_n731), .A3(new_n732), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n676), .A2(new_n366), .A3(new_n698), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n730), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n739), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n705), .A2(new_n708), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n813), .A4(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n919), .B(new_n920), .C1(new_n926), .C2(G953), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n369), .A2(new_n375), .ZN(new_n928));
  OR4_X1    g742(.A1(new_n928), .A2(new_n642), .A3(new_n736), .A4(new_n784), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n733), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n658), .A2(new_n813), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n924), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT126), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n930), .B(KEYINPUT125), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n936), .A2(new_n924), .A3(new_n938), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(G953), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n927), .B1(new_n945), .B2(new_n919), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n927), .C1(new_n945), .C2(new_n919), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  INV_X1    g767(.A(new_n913), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n926), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n289), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n287), .A2(new_n288), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n194), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n298), .B2(new_n299), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n808), .A2(new_n816), .A3(new_n953), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n861), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n940), .A2(new_n944), .A3(new_n913), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n962), .A2(new_n953), .B1(new_n288), .B2(new_n287), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n645), .ZN(G57));
endmodule


