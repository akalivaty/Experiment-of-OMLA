

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U324 ( .A1(n380), .A2(n580), .ZN(n382) );
  NAND2_X1 U325 ( .A1(n568), .A2(n435), .ZN(n436) );
  INV_X1 U326 ( .A(KEYINPUT112), .ZN(n381) );
  XNOR2_X1 U327 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U328 ( .A(n358), .B(n449), .ZN(n359) );
  XNOR2_X1 U329 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U330 ( .A(n392), .B(KEYINPUT48), .ZN(n545) );
  INV_X1 U331 ( .A(G169GAT), .ZN(n453) );
  XOR2_X1 U332 ( .A(n310), .B(n327), .Z(n572) );
  XNOR2_X1 U333 ( .A(n453), .B(KEYINPUT122), .ZN(n454) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n293) );
  XNOR2_X1 U336 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U338 ( .A(G113GAT), .B(G15GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G36GAT), .B(G50GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(G1GAT), .B(G8GAT), .Z(n297) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G197GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U345 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XOR2_X1 U346 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n301) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n424), .B(n302), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U352 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT70), .B(n309), .Z(n327) );
  XOR2_X1 U356 ( .A(KEYINPUT88), .B(G218GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(n313), .ZN(n433) );
  XOR2_X1 U360 ( .A(G8GAT), .B(G183GAT), .Z(n366) );
  XNOR2_X1 U361 ( .A(n433), .B(n366), .ZN(n315) );
  NAND2_X1 U362 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n318) );
  XOR2_X1 U364 ( .A(G64GAT), .B(G92GAT), .Z(n317) );
  XNOR2_X1 U365 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n357) );
  XOR2_X1 U367 ( .A(n318), .B(n357), .Z(n326) );
  XOR2_X1 U368 ( .A(KEYINPUT84), .B(KEYINPUT18), .Z(n320) );
  XNOR2_X1 U369 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U371 ( .A(n321), .B(KEYINPUT17), .Z(n323) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n323), .B(n322), .ZN(n443) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n324), .B(KEYINPUT77), .ZN(n337) );
  XNOR2_X1 U376 ( .A(n443), .B(n337), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n519) );
  INV_X1 U378 ( .A(n327), .ZN(n345) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT65), .B(KEYINPUT78), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U382 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n331) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(KEYINPUT66), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U385 ( .A(n333), .B(n332), .Z(n343) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(G85GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(KEYINPUT74), .ZN(n346) );
  XOR2_X1 U388 ( .A(n346), .B(G92GAT), .Z(n336) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U391 ( .A(n337), .B(G106GAT), .Z(n339) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(n418), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n345), .B(n344), .Z(n472) );
  XNOR2_X1 U398 ( .A(n346), .B(KEYINPUT72), .ZN(n348) );
  AND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U401 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n350) );
  XNOR2_X1 U402 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  NAND2_X1 U404 ( .A1(n352), .A2(n351), .ZN(n354) );
  OR2_X1 U405 ( .A1(n352), .A2(n351), .ZN(n353) );
  NAND2_X1 U406 ( .A1(n354), .A2(n353), .ZN(n360) );
  XOR2_X1 U407 ( .A(G78GAT), .B(G148GAT), .Z(n356) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n417) );
  XOR2_X1 U410 ( .A(n417), .B(n357), .Z(n358) );
  XOR2_X1 U411 ( .A(G120GAT), .B(G71GAT), .Z(n449) );
  XNOR2_X1 U412 ( .A(KEYINPUT13), .B(G57GAT), .ZN(n364) );
  XNOR2_X1 U413 ( .A(n361), .B(n364), .ZN(n577) );
  XNOR2_X1 U414 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n577), .B(n362), .ZN(n555) );
  NOR2_X1 U416 ( .A1(n555), .A2(n572), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n363), .B(KEYINPUT46), .ZN(n380) );
  XNOR2_X1 U418 ( .A(G71GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n379) );
  XOR2_X1 U420 ( .A(n366), .B(KEYINPUT79), .Z(n368) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U423 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n370) );
  XNOR2_X1 U424 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U427 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XOR2_X1 U428 ( .A(G64GAT), .B(G78GAT), .Z(n374) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(G155GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n448), .B(n375), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n559) );
  INV_X1 U434 ( .A(n559), .ZN(n580) );
  NOR2_X1 U435 ( .A1(n472), .A2(n383), .ZN(n384) );
  XNOR2_X1 U436 ( .A(KEYINPUT47), .B(n384), .ZN(n391) );
  XOR2_X1 U437 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n386) );
  INV_X1 U438 ( .A(n472), .ZN(n563) );
  XOR2_X1 U439 ( .A(KEYINPUT36), .B(n563), .Z(n583) );
  NAND2_X1 U440 ( .A1(n580), .A2(n583), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  NOR2_X1 U442 ( .A1(n387), .A2(n577), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n388), .B(KEYINPUT114), .ZN(n389) );
  NAND2_X1 U444 ( .A1(n389), .A2(n572), .ZN(n390) );
  NAND2_X1 U445 ( .A1(n391), .A2(n390), .ZN(n392) );
  NAND2_X1 U446 ( .A1(n519), .A2(n545), .ZN(n394) );
  XOR2_X1 U447 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n393) );
  XOR2_X1 U448 ( .A(n394), .B(n393), .Z(n568) );
  XOR2_X1 U449 ( .A(G155GAT), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT89), .B(KEYINPUT2), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n428) );
  XOR2_X1 U452 ( .A(G85GAT), .B(n428), .Z(n398) );
  NAND2_X1 U453 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U455 ( .A(G29GAT), .B(n399), .ZN(n416) );
  XOR2_X1 U456 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U459 ( .A(KEYINPUT92), .B(G57GAT), .Z(n403) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(G148GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U463 ( .A(G162GAT), .B(G127GAT), .Z(n407) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(G120GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U467 ( .A(n410), .B(KEYINPUT1), .Z(n414) );
  XOR2_X1 U468 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n412) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n446) );
  XNOR2_X1 U471 ( .A(n446), .B(KEYINPUT91), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n516) );
  INV_X1 U474 ( .A(n516), .ZN(n569) );
  XOR2_X1 U475 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n432) );
  XOR2_X1 U478 ( .A(G204GAT), .B(KEYINPUT22), .Z(n422) );
  XNOR2_X1 U479 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n423), .B(KEYINPUT85), .Z(n426) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT24), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U484 ( .A(n427), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U485 ( .A(n428), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n468) );
  AND2_X1 U489 ( .A1(n569), .A2(n468), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U491 ( .A(G176GAT), .B(G183GAT), .Z(n438) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n439), .B(KEYINPUT81), .Z(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(G190GAT), .Z(n441) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U502 ( .A(n451), .B(n450), .Z(n529) );
  INV_X1 U503 ( .A(n529), .ZN(n522) );
  NAND2_X1 U504 ( .A1(n452), .A2(n522), .ZN(n562) );
  NOR2_X1 U505 ( .A1(n572), .A2(n562), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n476) );
  NOR2_X1 U507 ( .A1(n572), .A2(n577), .ZN(n489) );
  XNOR2_X1 U508 ( .A(n519), .B(KEYINPUT94), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT27), .ZN(n466) );
  NOR2_X1 U510 ( .A1(n522), .A2(n468), .ZN(n458) );
  XNOR2_X1 U511 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n570) );
  NAND2_X1 U513 ( .A1(n466), .A2(n570), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n462) );
  NAND2_X1 U515 ( .A1(n522), .A2(n519), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT97), .B(n459), .Z(n460) );
  NAND2_X1 U517 ( .A1(n460), .A2(n468), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  AND2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n516), .A2(n465), .ZN(n471) );
  NAND2_X1 U521 ( .A1(n466), .A2(n516), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT95), .ZN(n543) );
  XOR2_X1 U523 ( .A(KEYINPUT28), .B(n468), .Z(n525) );
  INV_X1 U524 ( .A(n525), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n543), .A2(n469), .ZN(n528) );
  NOR2_X1 U526 ( .A1(n522), .A2(n528), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n486) );
  NOR2_X1 U528 ( .A1(n472), .A2(n559), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U530 ( .A1(n486), .A2(n474), .ZN(n503) );
  AND2_X1 U531 ( .A1(n489), .A2(n503), .ZN(n484) );
  NAND2_X1 U532 ( .A1(n484), .A2(n516), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U534 ( .A(n477), .B(KEYINPUT100), .Z(n479) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n484), .A2(n519), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT102), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U541 ( .A1(n484), .A2(n522), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n525), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT39), .Z(n492) );
  NOR2_X1 U546 ( .A1(n580), .A2(n486), .ZN(n487) );
  NAND2_X1 U547 ( .A1(n583), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n488), .ZN(n513) );
  NAND2_X1 U549 ( .A1(n513), .A2(n489), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n490), .Z(n498) );
  NAND2_X1 U551 ( .A1(n516), .A2(n498), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  XOR2_X1 U553 ( .A(G36GAT), .B(KEYINPUT103), .Z(n494) );
  NAND2_X1 U554 ( .A1(n519), .A2(n498), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n496) );
  NAND2_X1 U557 ( .A1(n522), .A2(n498), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n497), .Z(G1330GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U561 ( .A1(n498), .A2(n525), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n505) );
  INV_X1 U565 ( .A(n572), .ZN(n502) );
  NOR2_X1 U566 ( .A1(n502), .A2(n555), .ZN(n514) );
  AND2_X1 U567 ( .A1(n514), .A2(n503), .ZN(n509) );
  NAND2_X1 U568 ( .A1(n509), .A2(n516), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n519), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n522), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U576 ( .A1(n509), .A2(n525), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT109), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n524), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  XOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U585 ( .A1(n524), .A2(n519), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n545), .A2(n530), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n572), .A2(n539), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U597 ( .A1(n539), .A2(n555), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n559), .A2(n539), .ZN(n537) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n563), .A2(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  AND2_X1 U609 ( .A1(n570), .A2(n543), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n572), .A2(n553), .ZN(n546) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n555), .A2(n553), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n559), .A2(n553), .ZN(n552) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n563), .A2(n553), .ZN(n554) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n562), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n559), .A2(n562), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n567) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1351GAT) );
  AND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n576) );
  NOR2_X1 U637 ( .A1(n572), .A2(n576), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n576), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

