//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G119), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G119), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n192), .B2(new_n187), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(new_n189), .C1(new_n192), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT83), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT3), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(G104), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(new_n199), .A3(KEYINPUT83), .A4(G104), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G101), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(KEYINPUT84), .A3(G101), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  AND4_X1   g026(.A1(new_n212), .A2(new_n201), .A3(new_n203), .A4(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(new_n207), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n211), .A2(new_n215), .A3(KEYINPUT85), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT85), .B1(new_n211), .B2(new_n215), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n198), .B(new_n209), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT5), .B(new_n189), .C1(new_n192), .C2(new_n187), .ZN(new_n219));
  OR3_X1    g033(.A1(new_n188), .A2(KEYINPUT5), .A3(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(G113), .A3(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n201), .A2(new_n203), .A3(new_n212), .A4(new_n205), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n202), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n197), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n221), .A2(KEYINPUT89), .A3(new_n197), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(G110), .B(G122), .Z(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n218), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(KEYINPUT6), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n238), .A3(new_n233), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(KEYINPUT1), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n248));
  OAI221_X1 g062(.A(new_n243), .B1(G128), .B2(new_n244), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n244), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n245), .A2(G146), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n241), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n257), .B2(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n247), .A2(new_n259), .A3(new_n254), .A4(new_n255), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n251), .B1(new_n261), .B2(new_n250), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT90), .B(G224), .Z(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n262), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n237), .A2(new_n239), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(KEYINPUT7), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n270), .B(new_n271), .Z(new_n272));
  XOR2_X1   g086(.A(new_n233), .B(KEYINPUT8), .Z(new_n273));
  INV_X1    g087(.A(new_n227), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n226), .B1(new_n221), .B2(new_n197), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n236), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G210), .B1(G237), .B2(G902), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT92), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n267), .A2(new_n268), .A3(new_n279), .A4(new_n277), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n282), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT9), .B(G234), .Z(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(G217), .A3(new_n264), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n191), .A2(G122), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n188), .A2(G122), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G107), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n199), .A3(new_n291), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G128), .B(G143), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT13), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n242), .B2(G143), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n242), .A2(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT95), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n245), .A2(KEYINPUT13), .A3(G128), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(new_n306), .A3(KEYINPUT94), .A4(new_n301), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n304), .B2(new_n307), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n295), .B(new_n298), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT96), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n304), .A2(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT95), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n308), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT96), .A3(new_n298), .A4(new_n295), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n296), .B(new_n297), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n294), .B(KEYINPUT97), .Z(new_n320));
  INV_X1    g134(.A(KEYINPUT14), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n191), .A2(new_n321), .A3(G122), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT98), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n199), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n290), .A2(KEYINPUT14), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(KEYINPUT98), .A3(new_n291), .A4(new_n322), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT99), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT99), .B1(new_n324), .B2(new_n326), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n319), .B(new_n320), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n289), .B1(new_n318), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n329), .A3(new_n289), .ZN(new_n332));
  AOI21_X1  g146(.A(G902), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT100), .ZN(new_n334));
  INV_X1    g148(.A(G478), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT15), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n334), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n333), .B2(new_n334), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n264), .A2(G952), .ZN(new_n342));
  NAND2_X1  g156(.A1(G234), .A2(G237), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT21), .B(G898), .Z(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(G902), .A3(G953), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G475), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT16), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n250), .A3(G140), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n250), .A2(KEYINPUT16), .A3(G140), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT76), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n240), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(G146), .A3(new_n357), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n264), .A3(G214), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(new_n245), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT17), .A3(G131), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(G131), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n362), .B(G143), .ZN(new_n366));
  INV_X1    g180(.A(G131), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT17), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n359), .A2(new_n360), .A3(new_n364), .A4(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n351), .A2(KEYINPUT93), .A3(new_n353), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT93), .B1(new_n351), .B2(new_n353), .ZN(new_n373));
  OAI21_X1  g187(.A(G146), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n350), .B(KEYINPUT77), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n375), .A2(KEYINPUT78), .A3(new_n240), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT78), .B1(new_n375), .B2(new_n240), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(KEYINPUT18), .A2(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n363), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n223), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n371), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT19), .B1(new_n372), .B2(new_n373), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n240), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n365), .A2(new_n368), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n360), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n384), .B1(new_n382), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n348), .B(new_n268), .C1(new_n385), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT20), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n371), .A2(new_n382), .A3(new_n384), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n382), .A2(new_n391), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n348), .A4(new_n268), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n384), .B1(new_n371), .B2(new_n382), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n268), .B1(new_n385), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n394), .A2(new_n399), .B1(G475), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n341), .A2(new_n347), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G214), .B1(G237), .B2(G902), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT88), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n286), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G221), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n287), .B2(new_n268), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT82), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n268), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n264), .A2(G227), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n414), .B(new_n415), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n226), .B(new_n249), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT11), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n297), .B2(G137), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n297), .A2(G137), .ZN(new_n420));
  INV_X1    g234(.A(G137), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT11), .A3(G134), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G131), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n422), .A3(new_n367), .A4(new_n420), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT66), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n427), .A3(G131), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT12), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n226), .A2(new_n249), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n207), .A2(new_n214), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT4), .A3(new_n210), .A4(new_n222), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n211), .A2(new_n215), .A3(KEYINPUT85), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n208), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n261), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n435), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n429), .B(KEYINPUT86), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n416), .B1(new_n432), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT87), .B1(new_n443), .B2(new_n429), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n209), .B(new_n442), .C1(new_n216), .C2(new_n217), .ZN(new_n448));
  INV_X1    g262(.A(new_n435), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n430), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n416), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n443), .B2(new_n444), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n446), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n413), .B1(new_n456), .B2(G469), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n416), .B1(new_n453), .B2(new_n445), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(new_n432), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n412), .B(new_n268), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n411), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n426), .A2(new_n258), .A3(new_n260), .A4(new_n428), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n421), .A2(G134), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n420), .A3(KEYINPUT67), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n421), .A3(G134), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(G131), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT68), .A4(G131), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n249), .A2(new_n470), .A3(new_n425), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n472), .A3(KEYINPUT30), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n258), .B2(new_n260), .ZN(new_n476));
  XNOR2_X1  g290(.A(G143), .B(G146), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT0), .B(G128), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT64), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n253), .ZN(new_n480));
  AND4_X1   g294(.A1(new_n475), .A2(new_n479), .A3(new_n480), .A4(new_n260), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n474), .B1(new_n482), .B2(new_n430), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n198), .B(new_n473), .C1(new_n483), .C2(KEYINPUT30), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n463), .A2(new_n472), .A3(new_n197), .A4(new_n195), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(G101), .ZN(new_n487));
  INV_X1    g301(.A(G210), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n488), .A2(G237), .A3(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT31), .ZN(new_n493));
  INV_X1    g307(.A(new_n198), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n472), .A4(new_n463), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n485), .A2(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n494), .B2(new_n483), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n490), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT31), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n484), .A2(new_n501), .A3(new_n485), .A4(new_n491), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G472), .A2(G902), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT71), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n462), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n484), .A2(new_n508), .A3(new_n485), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n490), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n463), .A2(new_n472), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n198), .ZN(new_n513));
  INV_X1    g327(.A(new_n485), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n498), .A2(new_n513), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n516));
  INV_X1    g330(.A(G472), .ZN(new_n517));
  INV_X1    g331(.A(new_n481), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n430), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n472), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n496), .A2(new_n497), .B1(new_n521), .B2(new_n198), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n490), .A2(KEYINPUT29), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n510), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n517), .A2(new_n268), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n526), .B1(new_n525), .B2(new_n528), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n503), .A2(KEYINPUT32), .A3(new_n504), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n507), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(G119), .B2(new_n242), .ZN(new_n535));
  INV_X1    g349(.A(G119), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(KEYINPUT23), .A3(G128), .ZN(new_n537));
  OAI22_X1  g351(.A1(new_n535), .A2(new_n537), .B1(G119), .B2(new_n242), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G110), .ZN(new_n539));
  XOR2_X1   g353(.A(G119), .B(G128), .Z(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT74), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT24), .B(G110), .Z(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n356), .A2(G146), .A3(new_n357), .ZN(new_n544));
  AOI21_X1  g358(.A(G146), .B1(new_n356), .B2(new_n357), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n539), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n541), .A2(new_n542), .B1(G110), .B2(new_n538), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n360), .B(new_n547), .C1(new_n377), .C2(new_n376), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT22), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(G137), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n548), .A3(new_n552), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n268), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT25), .ZN(new_n557));
  INV_X1    g371(.A(G217), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(G234), .B2(new_n268), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n554), .A2(new_n560), .A3(new_n268), .A4(new_n555), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n565));
  INV_X1    g379(.A(new_n555), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n552), .B1(new_n546), .B2(new_n548), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n559), .A2(G902), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND4_X1   g384(.A1(new_n565), .A2(new_n554), .A3(new_n555), .A4(new_n569), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n557), .A2(KEYINPUT79), .A3(new_n559), .A4(new_n561), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n533), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(KEYINPUT81), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n533), .B2(new_n575), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n407), .B(new_n461), .C1(new_n577), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  OR2_X1    g395(.A1(new_n505), .A2(new_n506), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n503), .A2(new_n268), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n503), .A2(KEYINPUT101), .A3(new_n268), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(G472), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n461), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n574), .ZN(new_n589));
  INV_X1    g403(.A(new_n404), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n281), .B2(new_n283), .ZN(new_n591));
  INV_X1    g405(.A(new_n332), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT33), .B1(new_n592), .B2(new_n330), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n331), .A2(new_n594), .A3(new_n332), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n595), .A3(G478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n333), .A2(new_n335), .ZN(new_n597));
  NAND2_X1  g411(.A1(G478), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n402), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n591), .A2(new_n347), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n589), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  NAND2_X1  g418(.A1(new_n340), .A2(new_n339), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n337), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n393), .A2(KEYINPUT20), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT102), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n401), .A2(G475), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n394), .A2(new_n399), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n591), .A2(new_n347), .A3(new_n606), .A4(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT103), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT103), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n589), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  AND3_X1   g433(.A1(new_n341), .A2(new_n347), .A3(new_n402), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(new_n285), .A3(new_n284), .A4(new_n405), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n549), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n569), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n564), .A2(new_n573), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n621), .A2(new_n588), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT37), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G110), .ZN(G12));
  AND2_X1   g444(.A1(new_n591), .A2(new_n626), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n346), .A2(G900), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n344), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n608), .A2(new_n611), .A3(new_n609), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n341), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n631), .A2(new_n533), .A3(new_n461), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  INV_X1    g451(.A(new_n286), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n639), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n286), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n402), .B1(new_n605), .B2(new_n337), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n484), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n491), .B1(new_n645), .B2(new_n514), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n514), .B2(new_n511), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n513), .A2(new_n485), .A3(new_n490), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G472), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n507), .A2(new_n532), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n404), .A3(new_n627), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT106), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n286), .B(new_n639), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n655));
  INV_X1    g469(.A(new_n652), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .A4(new_n643), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n633), .B(KEYINPUT39), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n461), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT40), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n653), .A2(new_n657), .A3(KEYINPUT107), .A4(new_n661), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n245), .ZN(G45));
  AND2_X1   g481(.A1(new_n533), .A2(new_n461), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n669));
  INV_X1    g483(.A(new_n633), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n599), .A2(new_n402), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(new_n669), .A3(new_n631), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n533), .A2(new_n461), .A3(new_n591), .A4(new_n626), .ZN(new_n673));
  INV_X1    g487(.A(new_n671), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT108), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AND2_X1   g491(.A1(new_n533), .A2(new_n575), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n268), .B1(new_n458), .B2(new_n459), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n681));
  INV_X1    g495(.A(new_n409), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .A4(new_n460), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n680), .A2(new_n682), .A3(new_n460), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT109), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n678), .A2(new_n601), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n683), .A3(new_n685), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n614), .B2(new_n615), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n188), .ZN(G18));
  NAND2_X1  g505(.A1(new_n631), .A2(new_n533), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n685), .A2(new_n683), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n403), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n536), .ZN(G21));
  NAND2_X1  g509(.A1(new_n281), .A2(new_n283), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n404), .A3(new_n643), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n591), .A2(KEYINPUT111), .A3(new_n643), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n574), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n564), .A2(new_n572), .A3(KEYINPUT110), .A4(new_n573), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n515), .A2(new_n490), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n493), .A2(new_n706), .A3(new_n502), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n583), .A2(G472), .B1(new_n504), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n685), .A2(new_n347), .A3(new_n683), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT112), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  AND3_X1   g529(.A1(new_n671), .A2(new_n626), .A3(new_n708), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n685), .A2(new_n716), .A3(new_n591), .A4(new_n683), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n286), .A2(new_n719), .A3(new_n404), .A4(new_n671), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n409), .B1(new_n457), .B2(new_n460), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n533), .A2(new_n575), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n503), .A2(new_n504), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n462), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n531), .A2(new_n532), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n703), .A3(new_n704), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT113), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n703), .A3(new_n729), .A4(new_n704), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n286), .A2(new_n404), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n674), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n721), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n723), .B1(new_n734), .B2(KEYINPUT42), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NOR4_X1   g550(.A1(new_n722), .A2(new_n732), .A3(new_n341), .A4(new_n634), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n297), .ZN(G36));
  INV_X1    g552(.A(new_n399), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n609), .B1(new_n607), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n599), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT43), .Z(new_n742));
  AND2_X1   g556(.A1(new_n582), .A2(new_n587), .ZN(new_n743));
  OR3_X1    g557(.A1(new_n742), .A2(new_n743), .A3(new_n627), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n732), .A2(new_n658), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n453), .A2(new_n455), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n446), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(G469), .ZN(new_n752));
  INV_X1    g566(.A(new_n413), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n460), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n682), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n744), .A2(new_n745), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n746), .A2(new_n747), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(KEYINPUT114), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(KEYINPUT114), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n759), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(KEYINPUT114), .B(new_n764), .C1(new_n758), .C2(new_n682), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n533), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n574), .A4(new_n733), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NAND2_X1  g586(.A1(new_n680), .A2(new_n460), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n741), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n775), .A2(new_n776), .A3(new_n411), .A4(new_n705), .ZN(new_n777));
  INV_X1    g591(.A(new_n654), .ZN(new_n778));
  INV_X1    g592(.A(new_n651), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n405), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n742), .A2(new_n344), .A3(new_n705), .A4(new_n709), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n683), .A3(new_n685), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n590), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n732), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n781), .A2(KEYINPUT121), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT121), .B1(new_n781), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n773), .A2(new_n410), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n769), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n693), .A2(new_n732), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n574), .A2(new_n344), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n779), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n402), .A3(new_n599), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT122), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n799), .A3(new_n402), .A4(new_n599), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n742), .A2(new_n344), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n794), .A2(new_n802), .A3(new_n626), .A4(new_n708), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n787), .A2(new_n793), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n769), .A2(new_n792), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n807), .A2(new_n791), .B1(new_n785), .B2(new_n786), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n803), .A4(new_n801), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n806), .A2(new_n809), .A3(new_n342), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n781), .A2(new_n591), .A3(new_n683), .A4(new_n685), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n636), .A2(new_n717), .ZN(new_n812));
  AND4_X1   g626(.A1(KEYINPUT111), .A2(new_n696), .A3(new_n404), .A4(new_n643), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT111), .B1(new_n591), .B2(new_n643), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n651), .A2(new_n627), .A3(new_n633), .A4(new_n721), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n817), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT118), .B1(new_n819), .B2(new_n701), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n676), .B(new_n812), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(KEYINPUT120), .A3(new_n822), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n636), .A2(new_n717), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n820), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n819), .A2(new_n701), .A3(KEYINPUT118), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n676), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n286), .A2(new_n406), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n341), .B2(new_n740), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n606), .A2(KEYINPUT115), .A3(new_n402), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n743), .A2(new_n347), .A3(new_n575), .A4(new_n461), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n837), .B1(new_n845), .B2(new_n628), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n407), .A2(new_n461), .A3(new_n743), .A4(new_n626), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(KEYINPUT116), .C1(new_n844), .C2(new_n843), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n589), .A2(new_n838), .A3(new_n347), .A4(new_n600), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n580), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n854));
  INV_X1    g668(.A(new_n723), .ZN(new_n855));
  INV_X1    g669(.A(new_n737), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n634), .A2(new_n606), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n668), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n721), .A2(new_n671), .A3(new_n708), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n626), .A3(new_n788), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n694), .ZN(new_n863));
  INV_X1    g677(.A(new_n689), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n616), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n713), .A2(new_n863), .A3(new_n865), .A4(new_n686), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n853), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n836), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n821), .B(KEYINPUT52), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n723), .B(new_n737), .C1(new_n734), .C2(KEYINPUT42), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n851), .B1(new_n846), .B2(new_n848), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n686), .B1(new_n711), .B2(new_n712), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n690), .A3(new_n694), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n861), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n869), .B2(new_n874), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n810), .A2(new_n811), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n796), .A2(new_n600), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n794), .A2(new_n731), .A3(new_n802), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT48), .Z(new_n885));
  NOR3_X1   g699(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n780), .B1(new_n886), .B2(new_n887), .ZN(G75));
  AND2_X1   g702(.A1(new_n237), .A2(new_n239), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT123), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n266), .B(KEYINPUT55), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n268), .B1(new_n878), .B2(new_n879), .ZN(new_n894));
  AOI211_X1 g708(.A(KEYINPUT56), .B(new_n893), .C1(new_n894), .C2(G210), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n878), .A2(new_n879), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G210), .A3(G902), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n891), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n264), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n488), .B(new_n268), .C1(new_n878), .C2(new_n879), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n893), .B1(new_n903), .B2(KEYINPUT56), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n898), .A3(new_n892), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n890), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(G51));
  NAND2_X1  g721(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n881), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n753), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n753), .A2(KEYINPUT57), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n911), .A2(new_n912), .B1(new_n458), .B2(new_n459), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n894), .A2(G469), .A3(new_n750), .A4(new_n751), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n397), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n901), .ZN(G60));
  NAND2_X1  g734(.A1(new_n593), .A2(new_n595), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n598), .B(KEYINPUT59), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n877), .B2(new_n881), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n902), .C1(new_n921), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n878), .B2(new_n879), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n624), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n902), .B1(new_n930), .B2(new_n568), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n931), .B(new_n902), .C1(new_n568), .C2(new_n930), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT61), .B1(new_n936), .B2(KEYINPUT124), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(G66));
  AOI21_X1  g752(.A(new_n264), .B1(new_n263), .B2(new_n345), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n853), .A2(new_n866), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n264), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n891), .B1(G898), .B2(new_n264), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  NAND2_X1  g758(.A1(new_n771), .A2(new_n762), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n828), .A2(new_n830), .B1(new_n672), .B2(new_n675), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n664), .A2(new_n946), .A3(new_n665), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n664), .A2(new_n946), .A3(KEYINPUT62), .A4(new_n665), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n577), .A2(new_n579), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n842), .A2(new_n600), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n660), .A3(new_n788), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(G953), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n473), .B1(new_n483), .B2(KEYINPUT30), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT125), .Z(new_n957));
  AND2_X1   g771(.A1(new_n386), .A2(new_n388), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT126), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(G900), .A2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n945), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n760), .A2(new_n659), .A3(new_n701), .A4(new_n731), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n870), .A3(new_n946), .A4(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n960), .B(new_n962), .C1(new_n965), .C2(G953), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  INV_X1    g781(.A(new_n954), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n968), .B(new_n945), .C1(new_n949), .C2(new_n950), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n967), .B(new_n959), .C1(new_n969), .C2(G953), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n961), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT127), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G72));
  XNOR2_X1  g788(.A(new_n527), .B(KEYINPUT63), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n965), .B2(new_n941), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n645), .A2(new_n514), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n490), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n901), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n868), .A2(new_n876), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n646), .A3(new_n975), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n969), .A2(new_n940), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n646), .B1(new_n984), .B2(new_n975), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G57));
endmodule


