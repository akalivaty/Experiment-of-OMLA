//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n201), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G50), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n210), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n223), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G222), .A2(G1698), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT68), .B(G223), .Z(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n249), .A3(G274), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n249), .A2(new_n261), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT67), .B(G226), .Z(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G190), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(G200), .B2(new_n266), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n221), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n204), .A2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n210), .A2(G33), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT69), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n272), .B1(new_n279), .B2(KEYINPUT70), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(KEYINPUT70), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n271), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n210), .A3(G1), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n271), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n209), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n284), .B2(new_n271), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  MUX2_X1   g0091(.A(new_n285), .B(new_n291), .S(G50), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n282), .B2(new_n292), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n269), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n269), .C1(new_n294), .C2(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n293), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n266), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G179), .B2(new_n266), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n255), .B1(new_n209), .B2(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n286), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G77), .B2(new_n285), .ZN(new_n310));
  INV_X1    g0110(.A(new_n275), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n273), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n314), .B2(new_n271), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT3), .B(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G232), .A2(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G238), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G107), .C2(new_n316), .ZN(new_n322));
  INV_X1    g0122(.A(new_n264), .ZN(new_n323));
  INV_X1    g0123(.A(G274), .ZN(new_n324));
  INV_X1    g0124(.A(new_n221), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n248), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n323), .A2(G244), .B1(new_n326), .B2(new_n262), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n315), .B1(new_n303), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n322), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n315), .B(new_n333), .C1(new_n267), .C2(new_n328), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n307), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n311), .A2(new_n284), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n291), .B2(new_n311), .ZN(new_n337));
  INV_X1    g0137(.A(new_n271), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n341), .B2(new_n201), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n277), .A2(G159), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n316), .B2(G20), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(G68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n338), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n252), .A2(KEYINPUT73), .A3(G33), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n251), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n345), .A2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n340), .B1(new_n357), .B2(new_n346), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n351), .B1(new_n358), .B2(new_n344), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n337), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G232), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n263), .B1(new_n361), .B2(new_n264), .ZN(new_n362));
  OR2_X1    g0162(.A1(G223), .A2(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G226), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G1698), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n251), .A2(new_n363), .A3(new_n253), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n249), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n362), .A2(new_n368), .A3(new_n330), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n323), .A2(G232), .B1(new_n326), .B2(new_n262), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n321), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT18), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n316), .A2(new_n345), .A3(G20), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n254), .B2(new_n210), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n344), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n359), .A2(new_n380), .A3(new_n271), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n370), .B2(new_n372), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT74), .B(G190), .Z(new_n384));
  NOR3_X1   g0184(.A1(new_n362), .A2(new_n368), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n337), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n381), .A2(new_n387), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n373), .A2(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n330), .B2(new_n373), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n386), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n375), .A2(new_n390), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n286), .A2(G68), .A3(new_n288), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT72), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n340), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n274), .B2(new_n255), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n271), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n284), .A2(new_n340), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT12), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(KEYINPUT11), .A3(new_n271), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n400), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n263), .B1(new_n264), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n361), .A2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n316), .B(new_n414), .C1(G226), .C2(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n412), .B(new_n413), .C1(new_n417), .C2(new_n249), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n249), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT13), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G169), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(G179), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n421), .B2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n409), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n421), .A2(new_n267), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n382), .B1(new_n418), .B2(new_n420), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n428), .A2(new_n409), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n301), .A2(new_n335), .A3(new_n398), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G264), .A2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G257), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n316), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n252), .A2(G33), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n439));
  OAI21_X1  g0239(.A(G303), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n437), .A2(new_n440), .A3(KEYINPUT80), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT80), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n321), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n326), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n249), .ZN(new_n451));
  INV_X1    g0251(.A(G270), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n447), .B(new_n455), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n443), .A2(KEYINPUT81), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n384), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n321), .C1(new_n441), .C2(new_n442), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n210), .C1(G33), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n271), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n285), .A2(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n250), .A2(G1), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n284), .A2(new_n271), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(G116), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n454), .A2(new_n456), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n475), .A2(new_n460), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n461), .B(new_n474), .C1(new_n477), .C2(new_n382), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n330), .B1(new_n469), .B2(new_n473), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(new_n475), .A3(new_n460), .A4(new_n476), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n457), .A2(KEYINPUT82), .A3(new_n460), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n474), .A2(new_n303), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n475), .A2(new_n476), .A3(new_n460), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n478), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT6), .A3(G97), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n463), .A2(new_n491), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n206), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(KEYINPUT6), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n357), .A2(new_n346), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n491), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n271), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n285), .A2(G97), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n472), .B2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n447), .B1(new_n451), .B2(new_n435), .ZN(new_n504));
  INV_X1    g0304(.A(G244), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n251), .A3(new_n253), .A4(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(new_n462), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n251), .A3(new_n253), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT75), .B1(new_n510), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n249), .B1(new_n514), .B2(KEYINPUT76), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT76), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n516), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  AOI211_X1 g0317(.A(G190), .B(new_n504), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(KEYINPUT76), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(new_n321), .A3(new_n517), .ZN(new_n520));
  INV_X1    g0320(.A(new_n504), .ZN(new_n521));
  AOI21_X1  g0321(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n503), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n326), .A2(new_n445), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n249), .B(G250), .C1(G1), .C2(new_n444), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n250), .A2(new_n465), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n410), .A2(G1698), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n316), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT77), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n316), .A2(new_n532), .A3(G244), .A4(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n526), .B1(new_n534), .B2(new_n321), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT78), .B1(new_n535), .B2(new_n330), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n330), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n316), .A2(new_n210), .A3(G68), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n210), .B1(new_n416), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(G87), .B2(new_n207), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n273), .B2(new_n463), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n271), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n313), .A2(new_n284), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n313), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n472), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n534), .A2(new_n321), .ZN(new_n551));
  INV_X1    g0351(.A(new_n526), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n548), .A2(new_n550), .B1(new_n553), .B2(new_n303), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(G200), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n472), .A2(G87), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n546), .A2(new_n547), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(G190), .B2(new_n535), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n539), .A2(new_n554), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n507), .A2(new_n508), .A3(new_n462), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n510), .A2(new_n511), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n511), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n321), .B1(new_n565), .B2(new_n516), .ZN(new_n566));
  INV_X1    g0366(.A(new_n517), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n521), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n303), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n520), .A2(new_n330), .A3(new_n521), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n502), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n523), .A2(new_n559), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n251), .A2(new_n253), .A3(new_n210), .A4(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n316), .A2(new_n575), .A3(new_n210), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n210), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n491), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(new_n529), .B2(new_n210), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n578), .B1(new_n577), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n271), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n285), .B2(G107), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n491), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n472), .B2(G107), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(G250), .A2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n435), .A2(G1698), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(G294), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n595), .A2(new_n254), .B1(new_n250), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n321), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n450), .A2(G264), .A3(new_n249), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n447), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT84), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n602), .A3(new_n447), .A4(new_n599), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n603), .A3(G169), .ZN(new_n604));
  INV_X1    g0404(.A(new_n447), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n321), .B1(new_n445), .B2(new_n446), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n597), .A2(new_n321), .B1(new_n606), .B2(G264), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G179), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n592), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(G190), .B1(new_n601), .B2(new_n603), .ZN(new_n612));
  INV_X1    g0412(.A(new_n600), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n585), .B(new_n589), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR4_X1   g0416(.A1(new_n433), .A2(new_n490), .A3(new_n572), .A4(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n427), .A2(new_n332), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n390), .A3(new_n396), .A4(new_n430), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n375), .A2(new_n395), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n306), .B1(new_n621), .B2(new_n301), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n523), .A2(new_n571), .A3(new_n615), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n551), .A2(KEYINPUT85), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n534), .A2(new_n625), .A3(new_n321), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n526), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT87), .B1(new_n627), .B2(new_n382), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n535), .A2(G190), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n557), .B(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n534), .A2(new_n625), .A3(new_n321), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n534), .B2(new_n321), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n552), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(G200), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n628), .A2(new_n629), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT86), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n627), .B2(G169), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n548), .A2(new_n550), .B1(new_n535), .B2(new_n330), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n634), .A2(KEYINPUT86), .A3(new_n303), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n609), .A2(new_n590), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n484), .B(new_n644), .C1(new_n489), .C2(new_n488), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n623), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n571), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n637), .A3(new_n642), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n558), .A2(new_n555), .ZN(new_n650));
  INV_X1    g0450(.A(new_n538), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n536), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n548), .A2(new_n550), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(G169), .B2(new_n535), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n655), .B2(new_n571), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n642), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n646), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n622), .B1(new_n433), .B2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n611), .A2(new_n615), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n592), .A2(new_n610), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n615), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n668), .B2(new_n670), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n611), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n666), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n667), .A2(new_n474), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n490), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n484), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n489), .A2(new_n488), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT90), .B(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n667), .B1(new_n681), .B2(new_n682), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n672), .B2(new_n674), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n609), .A2(new_n590), .A3(new_n667), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n688), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n213), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n219), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n504), .B1(new_n515), .B2(new_n517), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT92), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n553), .A2(new_n608), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n477), .A2(new_n702), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n613), .A2(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n568), .A2(new_n708), .A3(new_n487), .A4(new_n634), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n535), .A2(G179), .A3(new_n607), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n487), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n705), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n666), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n706), .A2(new_n457), .A3(new_n460), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n704), .B1(new_n717), .B2(new_n568), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n709), .A3(new_n707), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n490), .A2(new_n572), .A3(new_n668), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n685), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n611), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n623), .A2(new_n643), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n642), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n655), .A2(new_n571), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n648), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n637), .A2(new_n642), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT26), .B1(new_n732), .B2(new_n571), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n623), .A2(new_n643), .A3(new_n725), .A4(KEYINPUT94), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n731), .B2(new_n733), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT29), .B(new_n667), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n667), .B1(new_n646), .B2(new_n657), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n724), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n701), .B1(new_n743), .B2(G1), .ZN(G364));
  XOR2_X1   g0544(.A(new_n687), .B(KEYINPUT95), .Z(new_n745));
  NOR2_X1   g0545(.A1(new_n283), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n209), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n696), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n745), .B(new_n750), .C1(new_n686), .C2(new_n684), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n695), .A2(new_n254), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G355), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G116), .B2(new_n213), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n695), .A2(new_n316), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n220), .B2(new_n444), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n243), .A2(new_n444), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n221), .B1(G20), .B2(new_n303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n749), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT98), .B1(new_n330), .B2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n210), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n330), .A2(KEYINPUT98), .A3(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n491), .ZN(new_n775));
  NAND2_X1  g0575(.A1(G20), .A2(G179), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n267), .A3(new_n382), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n775), .B1(G77), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n210), .B1(new_n784), .B2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n463), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(G20), .A3(new_n267), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OR3_X1    g0589(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT32), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n787), .A2(new_n790), .A3(new_n316), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n777), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(G68), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(new_n384), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n458), .A2(new_n382), .A3(new_n777), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n202), .B1(new_n339), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n770), .A2(new_n267), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G87), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n783), .A2(new_n795), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n774), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n788), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n316), .B1(new_n805), .B2(G329), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n596), .B2(new_n785), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(G322), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n778), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n796), .A2(G326), .B1(new_n810), .B2(G311), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n794), .A2(new_n812), .B1(new_n800), .B2(G303), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n802), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n766), .B1(new_n815), .B2(new_n763), .ZN(new_n816));
  INV_X1    g0616(.A(new_n762), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n684), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n751), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n334), .B1(new_n667), .B2(new_n315), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n332), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n332), .B2(new_n666), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n740), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n823), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n667), .B(new_n825), .C1(new_n646), .C2(new_n657), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n724), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n697), .B2(new_n747), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n724), .A2(new_n824), .A3(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n794), .A2(G283), .B1(new_n796), .B2(G303), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n781), .B2(new_n465), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT100), .Z(new_n833));
  INV_X1    g0633(.A(new_n774), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G87), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n316), .B(new_n786), .C1(G311), .C2(new_n805), .ZN(new_n837));
  INV_X1    g0637(.A(new_n800), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n491), .B2(new_n838), .C1(new_n596), .C2(new_n798), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n833), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n834), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n316), .B1(new_n788), .B2(new_n842), .C1(new_n339), .C2(new_n785), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n800), .B2(G50), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G143), .A2(new_n808), .B1(new_n796), .B2(G137), .ZN(new_n845));
  INV_X1    g0645(.A(new_n794), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n276), .B2(new_n846), .C1(new_n781), .C2(new_n789), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT34), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n841), .B(new_n844), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n763), .B1(new_n840), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n763), .A2(new_n760), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n750), .B1(new_n255), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(new_n761), .C2(new_n825), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n830), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n222), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  OR3_X1    g0660(.A1(new_n219), .A2(new_n255), .A3(new_n341), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n202), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n209), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n664), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n620), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n378), .A2(new_n379), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n351), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n337), .B1(new_n350), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n388), .B1(new_n870), .B2(new_n664), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n374), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n391), .A2(new_n394), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n391), .A2(new_n865), .ZN(new_n875));
  XNOR2_X1  g0675(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n388), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n870), .A2(new_n664), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n397), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n427), .A2(new_n666), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT105), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n874), .A2(new_n875), .A3(new_n388), .ZN(new_n887));
  INV_X1    g0687(.A(new_n876), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n664), .B1(new_n381), .B2(new_n387), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(KEYINPUT106), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n887), .A2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n397), .A2(new_n889), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n397), .A2(new_n896), .A3(new_n889), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n881), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n884), .B(new_n886), .C1(new_n900), .C2(KEYINPUT39), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n881), .A2(new_n882), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n409), .A2(new_n666), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n427), .A2(new_n430), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n427), .B2(new_n430), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n332), .A2(new_n666), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT101), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n826), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n902), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g0713(.A(KEYINPUT103), .B(new_n906), .C1(new_n826), .C2(new_n910), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n867), .B(new_n901), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n622), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n433), .B1(new_n740), .B2(new_n741), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n739), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n915), .B(new_n918), .Z(new_n919));
  INV_X1    g0719(.A(new_n903), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n431), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n427), .A2(new_n430), .A3(new_n903), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n823), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n721), .B2(new_n722), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n900), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n825), .B1(new_n904), .B2(new_n905), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT31), .B1(new_n719), .B2(new_n666), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n490), .ZN(new_n930));
  INV_X1    g0730(.A(new_n668), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n523), .A2(new_n559), .A3(new_n571), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n926), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n902), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n925), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n433), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n716), .A3(new_n720), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n937), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n686), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n919), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n209), .B2(new_n746), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n919), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n864), .B1(new_n944), .B2(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n691), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT109), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n503), .A2(new_n667), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n570), .A3(new_n569), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT108), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n523), .B(new_n571), .C1(new_n503), .C2(new_n667), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n948), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT109), .B1(new_n691), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n571), .B1(new_n957), .B2(new_n611), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(KEYINPUT42), .B1(new_n667), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT42), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n631), .A2(new_n667), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n643), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n642), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT43), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n964), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n688), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n957), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n961), .A2(new_n972), .A3(new_n971), .A4(new_n963), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT111), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n975), .A2(KEYINPUT111), .A3(new_n977), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n975), .A2(new_n978), .ZN(new_n984));
  INV_X1    g0784(.A(new_n977), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n981), .A2(new_n986), .A3(new_n987), .A4(new_n982), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n696), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n693), .B2(new_n957), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n692), .A4(new_n955), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT44), .B1(new_n693), .B2(new_n957), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n693), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n688), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n995), .B(new_n976), .C1(new_n996), .C2(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n675), .A2(new_n677), .A3(new_n689), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n691), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n687), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n745), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n743), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT112), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT112), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1000), .A4(new_n999), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n991), .B1(new_n1011), .B2(new_n743), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n989), .B(new_n990), .C1(new_n1012), .C2(new_n748), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n764), .B1(new_n213), .B2(new_n313), .C1(new_n756), .C2(new_n239), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(new_n749), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n771), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n846), .A2(new_n596), .B1(new_n1016), .B2(new_n463), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G311), .B2(new_n796), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n254), .B1(new_n788), .B2(new_n1019), .C1(new_n491), .C2(new_n785), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n808), .B2(G303), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n800), .A2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n782), .A2(G283), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(G143), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(new_n797), .B1(new_n846), .B2(new_n789), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G58), .B2(new_n800), .ZN(new_n1028));
  INV_X1    g0828(.A(G137), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n316), .B1(new_n788), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n771), .B2(G77), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1028), .B(new_n1031), .C1(new_n781), .C2(new_n202), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n785), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(G68), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n798), .B2(new_n276), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT113), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1025), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT47), .Z(new_n1038));
  INV_X1    g0838(.A(new_n763), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1015), .B1(new_n817), .B2(new_n968), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1013), .A2(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(G303), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n781), .A2(new_n1042), .B1(new_n1019), .B2(new_n798), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n794), .A2(G311), .B1(new_n796), .B2(G322), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n800), .A2(G294), .B1(G283), .B2(new_n1033), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT49), .Z(new_n1054));
  AOI21_X1  g0854(.A(new_n316), .B1(new_n805), .B2(G326), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1016), .B2(new_n465), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n785), .A2(new_n313), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n254), .B(new_n1058), .C1(G150), .C2(new_n805), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n789), .B2(new_n797), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n810), .A2(G68), .B1(new_n800), .B2(G77), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n202), .B2(new_n798), .C1(new_n275), .C2(new_n846), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(G97), .C2(new_n834), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n763), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n698), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n752), .A2(new_n1065), .B1(new_n491), .B2(new_n695), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n236), .A2(new_n444), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n311), .A2(new_n202), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n698), .B(new_n444), .C1(new_n340), .C2(new_n255), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n755), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1066), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n750), .B1(new_n1072), .B2(new_n764), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n678), .A2(new_n762), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n1075), .B1(new_n748), .B2(new_n1005), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1006), .A2(new_n696), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1005), .A2(new_n743), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  AOI21_X1  g0879(.A(new_n697), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1011), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n999), .A2(new_n748), .A3(new_n1000), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n755), .A2(new_n246), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n765), .B1(G97), .B2(new_n695), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n750), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G159), .A2(new_n808), .B1(new_n796), .B2(G150), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT51), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n311), .B2(new_n782), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n316), .B1(new_n788), .B2(new_n1026), .C1(new_n255), .C2(new_n785), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n800), .B2(G68), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n202), .B2(new_n846), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n836), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n316), .B1(new_n805), .B2(G322), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n465), .B2(new_n785), .C1(new_n838), .C2(new_n803), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n846), .A2(new_n1042), .B1(new_n596), .B2(new_n778), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n775), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G311), .A2(new_n808), .B1(new_n796), .B2(G317), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n1088), .A2(new_n1092), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1085), .B1(new_n1039), .B2(new_n1099), .C1(new_n955), .C2(new_n817), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1082), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1081), .A2(new_n1101), .ZN(G390));
  OAI21_X1  g0902(.A(new_n884), .B1(new_n900), .B2(KEYINPUT39), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n911), .B2(new_n886), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n667), .B(new_n825), .C1(new_n737), .C2(new_n738), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n906), .B1(new_n1105), .B2(new_n908), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n900), .A2(new_n886), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(G330), .B1(new_n721), .B2(new_n722), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(new_n926), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n906), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n724), .A2(new_n825), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1104), .B(new_n1113), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n748), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1103), .A2(new_n760), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n750), .B1(new_n275), .B2(new_n852), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n254), .B1(new_n788), .B2(new_n596), .C1(new_n255), .C2(new_n785), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G116), .A2(new_n808), .B1(new_n794), .B2(G107), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n803), .B2(new_n797), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G87), .C2(new_n800), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n841), .C1(new_n463), .C2(new_n781), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT120), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n254), .B1(new_n805), .B2(G125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n789), .B2(new_n785), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G128), .B2(new_n796), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n846), .A2(new_n1029), .B1(new_n1016), .B2(new_n202), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G132), .B2(new_n808), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n800), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT54), .B(G143), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n782), .A2(new_n1135), .ZN(new_n1136));
  AND4_X1   g0936(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1125), .A2(new_n1126), .A3(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1117), .B(new_n1118), .C1(new_n1039), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n724), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n906), .B1(new_n1142), .B2(new_n823), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1110), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(new_n1144), .B1(new_n826), .B2(new_n910), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(G330), .C1(new_n721), .C2(new_n722), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n825), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n939), .B2(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n906), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n908), .A3(new_n1105), .A4(new_n1113), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT117), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n723), .A2(new_n685), .A3(new_n906), .A4(new_n823), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1109), .A2(KEYINPUT116), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n825), .A3(new_n1148), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1155), .B1(new_n1157), .B2(new_n906), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1105), .A2(new_n908), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT117), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1146), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n739), .A2(new_n917), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n938), .A2(G330), .A3(new_n939), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n622), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n918), .A2(KEYINPUT115), .A3(new_n1163), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n697), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1161), .A2(new_n1168), .A3(new_n1114), .A4(new_n1111), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT118), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1158), .A2(KEYINPUT117), .A3(new_n1159), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1145), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1172), .A2(new_n1178), .A3(KEYINPUT118), .A4(new_n696), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1141), .B1(new_n1173), .B2(new_n1180), .ZN(G378));
  XOR2_X1   g0981(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n306), .B1(new_n298), .B2(new_n300), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n293), .A2(new_n865), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT55), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1183), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1182), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n937), .A2(G330), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n937), .B2(G330), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n915), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n935), .B1(new_n881), .B2(new_n882), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n924), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n896), .B1(new_n397), .B2(new_n889), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1201), .A2(new_n891), .A3(new_n892), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT38), .B1(new_n1202), .B2(new_n897), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n934), .B1(new_n1203), .B2(new_n881), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1200), .B1(new_n1204), .B2(KEYINPUT40), .ZN(new_n1205));
  INV_X1    g1005(.A(G330), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n826), .A2(new_n910), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1112), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT103), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n911), .A2(new_n912), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n902), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n901), .A2(new_n867), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n937), .A2(new_n1194), .A3(G330), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1207), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1197), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n748), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1189), .A2(new_n1192), .A3(new_n760), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n750), .B1(new_n202), .B2(new_n852), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1034), .B1(new_n797), .B2(new_n465), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT121), .Z(new_n1221));
  NOR2_X1   g1021(.A1(new_n316), .A2(G41), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n803), .B2(new_n788), .C1(new_n838), .C2(new_n255), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n808), .A2(G107), .B1(new_n771), .B2(G58), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n463), .B2(new_n846), .C1(new_n313), .C2(new_n778), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT122), .Z(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT58), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G33), .A2(G41), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1222), .A2(G50), .A3(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G128), .A2(new_n808), .B1(new_n796), .B2(G125), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n794), .A2(G132), .B1(new_n810), .B2(G137), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n800), .A2(new_n1135), .B1(G150), .B2(new_n1033), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n805), .A2(G124), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1230), .B(new_n1237), .C1(new_n1016), .C2(new_n789), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1235), .B2(KEYINPUT59), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1228), .A2(new_n1229), .A3(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1218), .B(new_n1219), .C1(new_n1241), .C2(new_n1039), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1217), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1177), .B1(new_n1115), .B2(new_n1161), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1197), .A2(new_n1215), .A3(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n915), .B(KEYINPUT125), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(KEYINPUT57), .A3(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n696), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1168), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1216), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n1250), .B2(new_n1252), .ZN(G375));
  AOI22_X1  g1053(.A1(new_n834), .A2(G77), .B1(new_n782), .B2(G107), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n254), .B1(new_n788), .B2(new_n1042), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1058), .B(new_n1255), .C1(new_n794), .C2(G116), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n797), .A2(new_n596), .B1(new_n803), .B2(new_n798), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G97), .B2(new_n800), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n797), .A2(new_n842), .B1(new_n1029), .B2(new_n798), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G159), .B2(new_n800), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n254), .B1(new_n805), .B2(G128), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n202), .B2(new_n785), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G58), .B2(new_n771), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n794), .A2(new_n1135), .B1(new_n810), .B2(G150), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1039), .B1(new_n1259), .B2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n750), .B(new_n1267), .C1(new_n340), .C2(new_n852), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1112), .B2(new_n761), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1176), .B2(new_n747), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(KEYINPUT126), .B(new_n1269), .C1(new_n1176), .C2(new_n747), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n991), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1169), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(G381));
  NAND3_X1  g1078(.A1(new_n1172), .A2(new_n1178), .A3(new_n696), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1141), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1076), .B(new_n819), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1281), .A2(G384), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(G381), .A2(new_n1280), .A3(G390), .A4(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1247), .A2(KEYINPUT57), .A3(new_n1248), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n697), .B1(new_n1284), .B2(new_n1251), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1251), .A2(new_n1216), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT57), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1243), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1283), .A2(new_n1040), .A3(new_n1013), .A4(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(new_n1280), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n665), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  AND3_X1   g1093(.A1(new_n1251), .A2(new_n1216), .A3(new_n1275), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1242), .B1(new_n1295), .B2(new_n747), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1141), .B(new_n1279), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT118), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1279), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1140), .B1(new_n1299), .B2(new_n1179), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1297), .B1(new_n1300), .B2(G375), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT60), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1276), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1176), .A2(KEYINPUT60), .A3(new_n1177), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n696), .A3(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1305), .A2(G384), .A3(new_n1274), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1305), .B2(new_n1274), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G213), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(G343), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1301), .A2(new_n1308), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1305), .A2(new_n1274), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n855), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1305), .A2(G384), .A3(new_n1274), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(G2897), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n1242), .B1(new_n747), .B2(new_n1295), .C1(new_n1286), .C2(new_n991), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(G378), .A2(new_n1289), .B1(new_n1291), .B2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1318), .B(new_n1320), .C1(new_n1322), .C2(new_n1310), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1301), .A2(new_n1308), .A3(new_n1325), .A4(new_n1311), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1313), .A2(new_n1323), .A3(new_n1324), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G393), .A2(G396), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(G390), .A2(new_n1281), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1281), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(new_n1081), .A3(new_n1101), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G387), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1013), .A2(new_n1329), .A3(new_n1040), .A4(new_n1331), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1327), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1335), .B1(new_n1337), .B2(new_n1312), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1320), .A2(new_n1318), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1301), .A2(new_n1311), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1312), .A2(new_n1337), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1338), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(new_n1343), .ZN(G405));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1333), .A2(new_n1345), .A3(new_n1334), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G378), .A2(new_n1289), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1291), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1308), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1347), .B(new_n1348), .C1(new_n1307), .C2(new_n1306), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1346), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1345), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1352), .B(new_n1353), .ZN(G402));
endmodule


