//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893;
  AND2_X1   g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n208), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n213), .A3(KEYINPUT71), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT66), .B(G183gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n221), .B1(new_n225), .B2(new_n222), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n228), .B(new_n229), .C1(new_n220), .C2(new_n223), .ZN(new_n230));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n232), .B1(KEYINPUT26), .B2(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n227), .A2(new_n230), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT24), .B1(new_n240), .B2(new_n222), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G190gat), .B2(new_n219), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n231), .B(KEYINPUT65), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n248), .A2(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(KEYINPUT64), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n231), .A4(new_n247), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n241), .A2(new_n243), .B1(new_n240), .B2(new_n222), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n256), .B2(KEYINPUT25), .ZN(new_n257));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n239), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n239), .A2(new_n257), .B1(new_n260), .B2(new_n258), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n217), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n217), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n239), .A2(new_n257), .A3(new_n258), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n265), .A2(KEYINPUT72), .A3(new_n267), .A4(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  AOI21_X1  g076(.A(KEYINPUT30), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  AOI211_X1 g079(.A(new_n279), .B(new_n280), .C1(new_n270), .C2(new_n271), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n271), .A3(new_n280), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n278), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT35), .ZN(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  INV_X1    g087(.A(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G113gat), .B2(G120gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G127gat), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n288), .B(new_n296), .C1(new_n291), .C2(new_n293), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(G134gat), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G155gat), .B(G162gat), .Z(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT75), .B(G162gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n303), .B1(new_n307), .B2(G155gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(G155gat), .B(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n302), .A3(new_n304), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(G134gat), .B1(new_n295), .B2(new_n297), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n298), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n297), .ZN(new_n315));
  INV_X1    g114(.A(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n295), .A2(G134gat), .A3(new_n297), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n287), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n298), .A2(new_n313), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n322), .B(new_n306), .C1(new_n308), .C2(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n318), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n312), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n319), .B1(KEYINPUT4), .B2(new_n286), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT5), .B(new_n320), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n319), .A2(KEYINPUT4), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n332), .A2(new_n327), .A3(new_n325), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT6), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n330), .A2(new_n340), .A3(new_n334), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n330), .B2(new_n334), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT6), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT85), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n284), .A2(new_n285), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G22gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n209), .B2(new_n213), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(KEYINPUT3), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n355), .A2(new_n311), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n323), .A2(new_n260), .B1(new_n214), .B2(new_n216), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n214), .A2(new_n260), .A3(new_n216), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n312), .B1(new_n359), .B2(new_n322), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361));
  NOR4_X1   g160(.A1(new_n360), .A2(new_n357), .A3(new_n361), .A4(new_n353), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n322), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n311), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n323), .A2(new_n260), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n353), .B1(new_n365), .B2(new_n217), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT78), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n352), .B(new_n358), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n358), .B1(new_n362), .B2(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G22gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT31), .ZN(new_n374));
  INV_X1    g173(.A(G50gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n369), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(new_n372), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n368), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n376), .B(KEYINPUT77), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT79), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n384), .B(new_n381), .C1(new_n372), .C2(new_n368), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n379), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n263), .A2(new_n326), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n239), .A2(new_n257), .A3(new_n321), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n394), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n390), .A3(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n397), .B(KEYINPUT32), .C1(new_n399), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n406), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n395), .A3(new_n393), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n386), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n351), .A2(new_n410), .A3(KEYINPUT86), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n284), .A2(new_n285), .A3(new_n350), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n408), .B(new_n396), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n386), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n344), .A2(new_n346), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n284), .A3(new_n386), .A4(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n411), .A2(new_n416), .B1(KEYINPUT35), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n386), .A2(KEYINPUT81), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n281), .A2(new_n283), .ZN(new_n421));
  INV_X1    g220(.A(new_n278), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n379), .B(new_n424), .C1(new_n383), .C2(new_n385), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n427));
  AND2_X1   g226(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n409), .B(new_n407), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n414), .B2(new_n428), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(KEYINPUT82), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n343), .A2(new_n342), .B1(new_n346), .B2(KEYINPUT85), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n277), .B1(new_n272), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n262), .A2(new_n268), .A3(KEYINPUT84), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT38), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n272), .A2(new_n277), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n434), .A2(new_n442), .A3(new_n443), .A4(new_n349), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT38), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n270), .A2(KEYINPUT37), .A3(new_n271), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n287), .B1(new_n328), .B2(new_n331), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n314), .A2(new_n319), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n286), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n341), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n287), .B(new_n454), .C1(new_n328), .C2(new_n331), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n453), .A2(KEYINPUT40), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT40), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n345), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n282), .B1(new_n443), .B2(new_n279), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n278), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(new_n386), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n432), .A2(new_n433), .B1(new_n448), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n419), .B1(new_n431), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n466), .B(G8gat), .Z(new_n467));
  INV_X1    g266(.A(KEYINPUT16), .ZN(new_n468));
  AOI21_X1  g267(.A(G1gat), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n467), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT14), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n475), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n477));
  XOR2_X1   g276(.A(G43gat), .B(G50gat), .Z(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n476), .A2(new_n480), .B1(new_n478), .B2(new_n477), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n481), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n470), .B(new_n484), .Z(new_n485));
  NAND2_X1  g284(.A1(G229gat), .A2(G233gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT89), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT13), .Z(new_n488));
  OR2_X1    g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n491), .A3(new_n483), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n484), .B2(new_n470), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT90), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(new_n494), .A2(new_n487), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n494), .B2(new_n487), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT11), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(new_n233), .ZN(new_n503));
  INV_X1    g302(.A(G197gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT12), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n489), .A2(new_n498), .A3(new_n506), .A4(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n463), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G57gat), .B(G64gat), .Z(new_n513));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514));
  INV_X1    g313(.A(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G71gat), .B(G78gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G127gat), .B(G155gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n470), .B1(new_n521), .B2(new_n520), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n240), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G211gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542));
  AND2_X1   g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n544), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n484), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(KEYINPUT41), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n490), .A2(new_n492), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT95), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n549), .A2(KEYINPUT41), .ZN(new_n559));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT93), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT96), .B1(new_n558), .B2(new_n562), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n555), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT97), .B1(new_n552), .B2(new_n555), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n557), .B(new_n561), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n536), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n547), .B(new_n520), .Z(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT98), .ZN(new_n575));
  INV_X1    g374(.A(new_n573), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n547), .A2(new_n520), .A3(new_n577), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G176gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(G204gat), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n575), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n574), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(KEYINPUT99), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n585), .B1(new_n590), .B2(new_n584), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n571), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n512), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n417), .B(KEYINPUT100), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT101), .B(G1gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(G1324gat));
  INV_X1    g396(.A(new_n593), .ZN(new_n598));
  INV_X1    g397(.A(new_n284), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT16), .B(G8gat), .Z(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT42), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(G8gat), .B1(new_n593), .B2(new_n284), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(G1325gat));
  NAND2_X1  g407(.A1(new_n409), .A2(new_n407), .ZN(new_n609));
  OR3_X1    g408(.A1(new_n593), .A2(G15gat), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(G15gat), .B1(new_n593), .B2(new_n430), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(G1326gat));
  NAND2_X1  g411(.A1(new_n420), .A2(new_n425), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT103), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n593), .B2(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT43), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G22gat), .ZN(G1327gat));
  INV_X1    g422(.A(new_n536), .ZN(new_n624));
  INV_X1    g423(.A(new_n591), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n510), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n432), .A2(new_n433), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n460), .B(new_n386), .C1(new_n444), .C2(new_n447), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n431), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n411), .A2(new_n416), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n418), .A2(KEYINPUT35), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n570), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT104), .B(KEYINPUT44), .C1(new_n463), .C2(new_n570), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n629), .A2(new_n426), .A3(new_n430), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n629), .A2(new_n426), .A3(KEYINPUT105), .A4(new_n430), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n633), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n569), .A2(new_n635), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n419), .B1(new_n641), .B2(new_n642), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n626), .B1(new_n638), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n594), .ZN(new_n654));
  INV_X1    g453(.A(new_n594), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n536), .A2(new_n570), .A3(new_n591), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n512), .A2(new_n471), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(G1328gat));
  OAI21_X1  g458(.A(G36gat), .B1(new_n653), .B2(new_n284), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n512), .A2(new_n472), .A3(new_n599), .A4(new_n656), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT46), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(G1329gat));
  INV_X1    g462(.A(G43gat), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n512), .A2(new_n664), .A3(new_n414), .A4(new_n656), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n653), .A2(new_n430), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(KEYINPUT47), .B(new_n665), .C1(new_n666), .C2(new_n664), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(G1330gat));
  INV_X1    g470(.A(KEYINPUT48), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n512), .A2(new_n375), .A3(new_n614), .A4(new_n656), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n375), .B1(new_n652), .B2(new_n614), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(KEYINPUT107), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n676), .B(new_n375), .C1(new_n652), .C2(new_n614), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n672), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G50gat), .B1(new_n653), .B2(new_n386), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT48), .A3(new_n673), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n511), .A2(new_n591), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n649), .A2(new_n571), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n655), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n599), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT49), .B(G64gat), .Z(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(G1333gat));
  NAND3_X1  g488(.A1(new_n683), .A2(new_n515), .A3(new_n414), .ZN(new_n690));
  INV_X1    g489(.A(new_n430), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n515), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n694), .A2(KEYINPUT50), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT50), .B1(new_n694), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(G1334gat));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n614), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g499(.A1(new_n536), .A2(new_n510), .A3(new_n570), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n644), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n644), .A2(KEYINPUT51), .A3(new_n701), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n625), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(G85gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n707), .A3(new_n655), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n638), .A2(new_n651), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n624), .A2(new_n511), .A3(new_n591), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n594), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n714), .B(new_n708), .C1(new_n711), .C2(new_n707), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1336gat));
  INV_X1    g515(.A(G92gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(new_n717), .A3(new_n599), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n709), .A2(new_n284), .A3(new_n710), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT52), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n718), .C1(new_n719), .C2(new_n717), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1337gat));
  XNOR2_X1  g523(.A(KEYINPUT110), .B(G99gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n414), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n430), .A3(new_n710), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT111), .B(new_n726), .C1(new_n727), .C2(new_n725), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1338gat));
  INV_X1    g531(.A(G106gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n386), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n706), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n709), .A2(new_n710), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n614), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(G106gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n733), .B1(new_n736), .B2(new_n734), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(G1339gat));
  NAND3_X1  g541(.A1(new_n578), .A2(new_n576), .A3(new_n579), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT54), .B(new_n581), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n587), .A2(new_n748), .A3(new_n589), .ZN(new_n749));
  INV_X1    g548(.A(new_n584), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n747), .A2(new_n749), .A3(KEYINPUT55), .A4(new_n750), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n753), .A2(new_n510), .A3(new_n585), .A4(new_n754), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n485), .A2(new_n488), .B1(new_n494), .B2(new_n487), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n756), .A2(KEYINPUT113), .A3(new_n505), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n756), .B2(new_n505), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(new_n509), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n591), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n569), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n569), .A2(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n753), .A2(new_n585), .A3(new_n754), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n624), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n536), .A2(new_n511), .A3(new_n570), .A4(new_n625), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n594), .A2(new_n599), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n609), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n768), .A2(new_n613), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G113gat), .B1(new_n774), .B2(new_n511), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n415), .A2(new_n599), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n768), .A2(new_n655), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n510), .A2(new_n289), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT115), .Z(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(G1340gat));
  NOR3_X1   g579(.A1(new_n774), .A2(new_n290), .A3(new_n625), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n777), .A2(new_n625), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n290), .B2(new_n782), .ZN(G1341gat));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n536), .A2(G127gat), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n774), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n296), .B1(new_n777), .B2(new_n624), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n774), .B2(new_n785), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT117), .ZN(G1342gat));
  OAI21_X1  g589(.A(G134gat), .B1(new_n774), .B2(new_n570), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n569), .A2(new_n316), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n777), .A2(KEYINPUT56), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT56), .B1(new_n777), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n791), .B(KEYINPUT118), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n796), .A4(new_n795), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1343gat));
  NOR3_X1   g601(.A1(new_n691), .A2(new_n386), .A3(new_n599), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n768), .A2(new_n655), .A3(new_n770), .A4(new_n803), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n804), .A2(G141gat), .A3(new_n511), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n768), .A2(new_n734), .A3(new_n770), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n765), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n765), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n766), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n613), .A2(new_n807), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n806), .A2(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n772), .A2(new_n691), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT120), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n813), .A2(new_n511), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n805), .B1(new_n817), .B2(new_n300), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n805), .B2(KEYINPUT122), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n805), .B1(KEYINPUT122), .B2(new_n819), .C1(new_n817), .C2(new_n300), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1344gat));
  OR4_X1    g622(.A1(KEYINPUT59), .A2(new_n813), .A3(new_n625), .A4(new_n816), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n613), .A2(KEYINPUT57), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n806), .A2(KEYINPUT57), .B1(new_n767), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n591), .A3(new_n815), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT59), .B1(new_n804), .B2(new_n625), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n301), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n828), .A3(new_n830), .ZN(G1345gat));
  NOR3_X1   g630(.A1(new_n813), .A2(new_n624), .A3(new_n816), .ZN(new_n832));
  INV_X1    g631(.A(G155gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n536), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n832), .A2(new_n833), .B1(new_n804), .B2(new_n834), .ZN(G1346gat));
  OR3_X1    g634(.A1(new_n804), .A2(new_n307), .A3(new_n570), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n813), .A2(new_n570), .A3(new_n816), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n307), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(G1347gat));
  NOR2_X1   g640(.A1(new_n655), .A2(new_n284), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n414), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n768), .A2(new_n613), .A3(new_n845), .A4(new_n770), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n233), .A3(new_n511), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n410), .A2(new_n768), .A3(new_n770), .A4(new_n842), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n510), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n233), .ZN(G1348gat));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n234), .A3(new_n591), .ZN(new_n851));
  OAI21_X1  g650(.A(G176gat), .B1(new_n846), .B2(new_n625), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1349gat));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n225), .A3(new_n536), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n219), .B1(new_n846), .B2(new_n624), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g656(.A(G190gat), .B1(new_n846), .B2(new_n570), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT125), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(G190gat), .C1(new_n846), .C2(new_n570), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(KEYINPUT61), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n848), .A2(new_n222), .A3(new_n569), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n858), .A2(KEYINPUT125), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n862), .A2(KEYINPUT126), .A3(new_n863), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1351gat));
  INV_X1    g669(.A(new_n842), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n691), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n806), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(G197gat), .B1(new_n874), .B2(new_n510), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n826), .A2(new_n872), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n511), .A2(new_n504), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1352gat));
  INV_X1    g677(.A(new_n874), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n625), .A2(G204gat), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT62), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT127), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n826), .A2(new_n591), .A3(new_n872), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G204gat), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n879), .A2(KEYINPUT62), .A3(new_n880), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(G1353gat));
  OR3_X1    g685(.A1(new_n879), .A2(G211gat), .A3(new_n624), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n826), .A2(new_n536), .A3(new_n872), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT63), .B1(new_n888), .B2(G211gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(G1354gat));
  AOI21_X1  g690(.A(G218gat), .B1(new_n874), .B2(new_n569), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n569), .A2(G218gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n876), .B2(new_n893), .ZN(G1355gat));
endmodule


