//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(G101), .B1(new_n192), .B2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n193), .A2(new_n200), .A3(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(new_n199), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n192), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n221), .B2(new_n198), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n201), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(G128), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G143), .B2(new_n209), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n213), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n210), .A3(new_n212), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n230), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n236), .B2(new_n207), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n201), .A4(new_n222), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n222), .A2(new_n201), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n241), .B2(new_n237), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n224), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT80), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n246), .A2(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n231), .A2(new_n210), .A3(new_n212), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT79), .B1(new_n249), .B2(new_n223), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n239), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT80), .A3(new_n224), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n235), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT11), .A3(G134), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G131), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT65), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n254), .A2(KEYINPUT11), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n258), .A2(new_n259), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n259), .B1(new_n258), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n253), .A2(KEYINPUT85), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n205), .A2(new_n219), .B1(new_n233), .B2(new_n225), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT80), .B1(new_n251), .B2(new_n224), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n244), .B(KEYINPUT10), .C1(new_n250), .C2(new_n239), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n268), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n268), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n245), .A2(new_n252), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT81), .A3(new_n268), .A4(new_n271), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G110), .B(G140), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT78), .ZN(new_n285));
  INV_X1    g099(.A(G227), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G953), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n285), .B(new_n287), .Z(new_n288));
  NOR3_X1   g102(.A1(new_n277), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n282), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n251), .B1(new_n241), .B2(new_n233), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n275), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT83), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n291), .A2(new_n295), .A3(new_n275), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n275), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT12), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n305), .B2(new_n288), .ZN(new_n306));
  OAI21_X1  g120(.A(G469), .B1(new_n306), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  INV_X1    g122(.A(new_n288), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT85), .B1(new_n253), .B2(new_n268), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n274), .A2(new_n270), .A3(new_n275), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(new_n290), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n290), .A2(new_n309), .A3(new_n300), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n308), .B(new_n190), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT86), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n290), .A2(new_n309), .A3(new_n300), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n310), .A2(new_n311), .B1(new_n280), .B2(new_n282), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n308), .A4(new_n190), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n191), .B1(new_n307), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n229), .A2(new_n325), .A3(new_n232), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT91), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT91), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n229), .A2(new_n328), .A3(new_n325), .A4(new_n232), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n218), .B2(G125), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n218), .A2(new_n332), .A3(G125), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI211_X1 g150(.A(KEYINPUT89), .B(new_n325), .C1(new_n208), .C2(new_n217), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n333), .A2(new_n337), .A3(KEYINPUT90), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(G224), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G224), .ZN(new_n342));
  OAI221_X1 g156(.A(new_n330), .B1(new_n342), .B2(G953), .C1(new_n336), .C2(new_n338), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G116), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT67), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G116), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(G119), .ZN(new_n349));
  INV_X1    g163(.A(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G116), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT2), .B(G113), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n351), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT68), .B1(new_n349), .B2(new_n351), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G113), .B1(new_n351), .B2(KEYINPUT5), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n241), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n355), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n205), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n352), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n351), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(KEYINPUT5), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n360), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n372), .A2(KEYINPUT87), .A3(new_n241), .A4(new_n355), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G122), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n363), .A2(new_n366), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n363), .A2(new_n366), .A3(new_n373), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AOI22_X1  g192(.A1(KEYINPUT6), .A2(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n366), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n354), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT87), .B1(new_n381), .B2(new_n241), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT6), .B(new_n378), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n344), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT7), .B1(new_n342), .B2(G953), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n330), .B(new_n387), .C1(new_n336), .C2(new_n338), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n330), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n333), .A2(new_n337), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n327), .A2(KEYINPUT92), .A3(new_n329), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n386), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n223), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n374), .B(KEYINPUT8), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n349), .A2(KEYINPUT5), .A3(new_n351), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n354), .B1(new_n371), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n395), .B(new_n396), .C1(new_n223), .C2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n375), .A2(new_n388), .A3(new_n394), .A4(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n400), .A2(new_n190), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n385), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n385), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n324), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n323), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n208), .B(new_n217), .C1(new_n266), .C2(new_n267), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n258), .A2(new_n259), .A3(new_n265), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n259), .B1(G134), .B2(G137), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n261), .A2(new_n263), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G137), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n233), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n408), .A2(new_n355), .A3(new_n364), .A4(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n416));
  NOR2_X1   g230(.A1(G237), .A2(G953), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G210), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT26), .B(G101), .Z(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n365), .ZN(new_n423));
  INV_X1    g237(.A(new_n267), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n218), .B1(new_n424), .B2(new_n409), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n233), .A2(new_n409), .A3(new_n412), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT30), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n408), .A2(new_n428), .A3(new_n413), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n423), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n414), .A2(new_n421), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT70), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT31), .ZN(new_n435));
  INV_X1    g249(.A(new_n421), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n365), .B1(new_n425), .B2(new_n426), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n414), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT28), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT28), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n414), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n437), .B2(new_n414), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n439), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n436), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n408), .A2(new_n428), .A3(new_n413), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n428), .B1(new_n408), .B2(new_n413), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n365), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT31), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n414), .A2(new_n421), .A3(new_n415), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n433), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n435), .B(new_n446), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(G472), .A2(G902), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(KEYINPUT32), .A3(new_n457), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n443), .A2(new_n445), .A3(new_n436), .ZN(new_n462));
  INV_X1    g276(.A(new_n414), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n436), .B1(new_n430), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n462), .A2(KEYINPUT29), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n442), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(new_n444), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n421), .A2(KEYINPUT29), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(KEYINPUT73), .A3(new_n469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n190), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G472), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n460), .A2(new_n461), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n417), .A2(G214), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n211), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n417), .A2(G143), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT18), .A2(G131), .ZN(new_n482));
  INV_X1    g296(.A(G140), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n325), .A2(G140), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G146), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(G146), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n481), .A2(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n481), .A2(new_n491), .A3(new_n482), .ZN(new_n492));
  INV_X1    g306(.A(new_n482), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT93), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT16), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n496), .A2(G146), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(G146), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n480), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n480), .A2(G131), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n478), .A2(new_n259), .A3(new_n479), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n500), .B(new_n501), .C1(new_n504), .C2(KEYINPUT17), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n192), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT95), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(KEYINPUT94), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n513), .A3(new_n503), .ZN(new_n514));
  XNOR2_X1  g328(.A(G125), .B(G140), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT19), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n498), .B1(new_n516), .B2(new_n209), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n507), .B1(new_n518), .B2(new_n495), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n511), .A2(new_n519), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n524), .B2(KEYINPUT96), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(KEYINPUT96), .A3(new_n523), .A4(new_n521), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n507), .B1(new_n495), .B2(new_n505), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n190), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(KEYINPUT97), .ZN(new_n531));
  INV_X1    g345(.A(G475), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n530), .B2(KEYINPUT97), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n346), .A2(new_n348), .A3(G122), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT99), .B1(new_n536), .B2(KEYINPUT14), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT98), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n345), .B2(G122), .ZN(new_n539));
  INV_X1    g353(.A(G122), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT98), .A3(G116), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n536), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g359(.A(G107), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n226), .A2(G143), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n211), .A2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n411), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n547), .A2(new_n261), .A3(new_n263), .A4(new_n548), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n542), .A2(new_n536), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n195), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n548), .B(KEYINPUT13), .Z(new_n555));
  INV_X1    g369(.A(new_n547), .ZN(new_n556));
  OAI21_X1  g370(.A(G134), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n552), .A2(new_n195), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n552), .A2(new_n195), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n551), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G217), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n188), .A2(new_n562), .A3(G953), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n560), .A3(new_n563), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n340), .A2(G952), .ZN(new_n573));
  NAND2_X1  g387(.A1(G234), .A2(G237), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(G902), .A3(G953), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n535), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n562), .B1(G234), .B2(new_n190), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT23), .B1(new_n230), .B2(G119), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT74), .B1(new_n350), .B2(G128), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n230), .A3(G119), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT66), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G128), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n590), .A3(KEYINPUT23), .A4(G119), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT76), .B(G110), .Z(new_n592));
  AND3_X1   g406(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT24), .B(G110), .Z(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(new_n590), .A3(G119), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n350), .A2(G128), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n515), .B2(KEYINPUT16), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G146), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n488), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT77), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n498), .A2(new_n487), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n604), .B(new_n605), .C1(new_n597), .C2(new_n593), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT75), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n498), .B2(new_n499), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n587), .A2(new_n591), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(G110), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n496), .A2(new_n497), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n209), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n601), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(G110), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(KEYINPUT75), .A3(new_n617), .A4(new_n609), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT22), .B(G137), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n620), .B(new_n621), .Z(new_n622));
  AND3_X1   g436(.A1(new_n607), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n607), .B2(new_n619), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT25), .B1(new_n625), .B2(new_n190), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NOR4_X1   g441(.A1(new_n623), .A2(new_n624), .A3(new_n627), .A4(G902), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n582), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n582), .A2(G902), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n476), .A2(new_n581), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n407), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n456), .A2(new_n190), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n456), .B2(new_n190), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n632), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n323), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n580), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n526), .A2(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n565), .A2(new_n566), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT33), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n565), .A2(new_n648), .A3(new_n566), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n649), .A3(G478), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n568), .A2(new_n190), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n567), .B2(new_n568), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n385), .A2(new_n401), .ZN(new_n655));
  INV_X1    g469(.A(new_n402), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n385), .A2(new_n401), .A3(new_n402), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT101), .B1(new_n659), .B2(new_n324), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  INV_X1    g475(.A(new_n324), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n661), .B(new_n662), .C1(new_n657), .C2(new_n658), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n644), .B(new_n654), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n643), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT34), .B(G104), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n522), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n522), .B1(new_n670), .B2(KEYINPUT20), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n669), .A2(new_n671), .B1(new_n570), .B2(new_n571), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n580), .B(KEYINPUT103), .Z(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n534), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n405), .A2(new_n661), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n324), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n643), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT35), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NAND2_X1  g495(.A1(new_n607), .A2(new_n619), .ZN(new_n682));
  INV_X1    g496(.A(new_n622), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n682), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n630), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n629), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n572), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n645), .A3(new_n644), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n641), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n407), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  OR2_X1    g507(.A1(new_n577), .A2(G900), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n575), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n531), .B2(new_n533), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n672), .A2(new_n687), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n675), .B2(new_n676), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n288), .B1(new_n277), .B2(new_n283), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n700), .B2(new_n317), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n320), .B1(new_n701), .B2(new_n308), .ZN(new_n702));
  INV_X1    g516(.A(new_n321), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n300), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT84), .B1(new_n290), .B2(new_n300), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n288), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n289), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI22_X1  g522(.A1(new_n702), .A2(new_n703), .B1(new_n708), .B2(new_n308), .ZN(new_n709));
  INV_X1    g523(.A(new_n191), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n699), .A2(new_n709), .A3(new_n710), .A4(new_n476), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT104), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n323), .A2(new_n713), .A3(new_n476), .A4(new_n699), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G128), .ZN(G30));
  XNOR2_X1  g530(.A(new_n695), .B(KEYINPUT39), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n323), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT40), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n718), .B(KEYINPUT40), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT106), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n659), .B(KEYINPUT38), .Z(new_n725));
  INV_X1    g539(.A(new_n461), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n456), .B2(new_n457), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n438), .A2(new_n436), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n434), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(G902), .B1(new_n730), .B2(KEYINPUT105), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(KEYINPUT105), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G472), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n645), .A2(new_n688), .ZN(new_n735));
  INV_X1    g549(.A(new_n687), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n324), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n725), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n722), .A2(new_n724), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  NOR3_X1   g554(.A1(new_n645), .A2(new_n653), .A3(new_n696), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n687), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n675), .B2(new_n676), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n323), .A2(new_n476), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT107), .B(G146), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G48));
  NAND2_X1  g560(.A1(new_n476), .A2(new_n633), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n308), .B1(new_n319), .B2(new_n190), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n191), .B(new_n749), .C1(new_n316), .C2(new_n321), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n654), .A2(new_n644), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n675), .B2(new_n676), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n749), .B1(new_n316), .B2(new_n321), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n710), .A3(new_n476), .A4(new_n633), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n678), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n748), .A2(new_n750), .A3(new_n677), .A4(KEYINPUT108), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  NAND2_X1  g576(.A1(new_n675), .A2(new_n676), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n757), .A3(new_n710), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n476), .A2(new_n581), .A3(new_n687), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT109), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n765), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n750), .A3(new_n768), .A4(new_n763), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  INV_X1    g585(.A(new_n735), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n675), .B2(new_n676), .ZN(new_n773));
  INV_X1    g587(.A(G472), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n456), .B2(new_n190), .ZN(new_n775));
  INV_X1    g589(.A(new_n457), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n431), .A2(KEYINPUT71), .A3(new_n450), .A4(new_n433), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n452), .A2(new_n453), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n778), .B1(new_n434), .B2(KEYINPUT31), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n436), .B1(new_n467), .B2(new_n444), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n673), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n775), .A2(new_n781), .A3(new_n632), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n750), .A2(new_n773), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G122), .ZN(G24));
  NOR2_X1   g599(.A1(new_n775), .A2(new_n781), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n687), .A3(new_n741), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n764), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n325), .ZN(G27));
  NAND3_X1  g603(.A1(new_n657), .A2(new_n324), .A3(new_n658), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n323), .A2(new_n748), .A3(new_n741), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n191), .B(new_n790), .C1(new_n307), .C2(new_n322), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT42), .A3(new_n748), .A4(new_n741), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n259), .ZN(G33));
  AND2_X1   g616(.A1(new_n672), .A2(new_n697), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n323), .A2(new_n748), .A3(new_n803), .A4(new_n791), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND2_X1  g619(.A1(new_n306), .A2(KEYINPUT45), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n309), .B1(new_n303), .B2(new_n304), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n289), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(G469), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(G469), .A2(G902), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n812), .A2(KEYINPUT46), .B1(new_n321), .B2(new_n316), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n812), .B2(KEYINPUT46), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n811), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(KEYINPUT111), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n790), .B(KEYINPUT113), .Z(new_n820));
  NOR3_X1   g634(.A1(new_n535), .A2(new_n653), .A3(KEYINPUT43), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n653), .B1(new_n535), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n645), .A2(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n825), .B2(KEYINPUT43), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n641), .A3(new_n687), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT44), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n829), .A3(new_n641), .A4(new_n687), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n820), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n819), .A2(new_n710), .A3(new_n717), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(KEYINPUT114), .B(G137), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(G39));
  NAND2_X1  g648(.A1(new_n819), .A2(new_n710), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n819), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n460), .A2(new_n461), .A3(new_n475), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n840), .A2(new_n632), .A3(new_n741), .A4(new_n791), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  INV_X1    g657(.A(new_n734), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n633), .A2(new_n710), .A3(new_n324), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n825), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n757), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n725), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n750), .A2(new_n576), .A3(new_n791), .A4(new_n826), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n748), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT48), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n632), .A2(new_n575), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n734), .A2(new_n750), .A3(new_n791), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n654), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n826), .A2(new_n576), .A3(new_n633), .A4(new_n786), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(new_n764), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n573), .A2(new_n854), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n687), .A3(new_n786), .ZN(new_n861));
  NAND2_X1  g675(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n725), .A2(new_n750), .A3(new_n662), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(new_n858), .ZN(new_n864));
  NOR2_X1   g678(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n645), .A2(new_n653), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n864), .A2(new_n865), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n861), .A2(KEYINPUT51), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n847), .A2(new_n710), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n837), .A2(new_n838), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n858), .A2(new_n820), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI211_X1 g690(.A(KEYINPUT120), .B(new_n869), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n838), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n871), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT116), .B1(new_n837), .B2(new_n838), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n861), .A2(new_n866), .A3(new_n868), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT119), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n788), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n715), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n788), .B1(new_n712), .B2(new_n714), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n736), .A2(new_n695), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n728), .B2(new_n733), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n323), .A2(new_n893), .A3(new_n773), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n744), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT52), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT52), .B1(new_n889), .B2(new_n895), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n323), .B(new_n406), .C1(new_n634), .C2(new_n690), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n654), .B1(new_n645), .B2(new_n572), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n405), .A3(new_n782), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n323), .A2(new_n904), .A3(new_n642), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n572), .B1(new_n669), .B2(new_n671), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n687), .A3(new_n697), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n787), .B1(new_n840), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n323), .A3(new_n791), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n804), .A2(new_n902), .A3(new_n905), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n749), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n783), .A2(new_n322), .A3(new_n710), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n735), .B1(new_n660), .B2(new_n663), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n758), .A2(new_n664), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n759), .B2(new_n760), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n910), .A2(new_n915), .A3(new_n770), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n801), .A2(new_n916), .A3(KEYINPUT53), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n901), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n895), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n899), .ZN(new_n920));
  INV_X1    g734(.A(new_n914), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n761), .A2(new_n770), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n799), .A3(new_n800), .A4(new_n910), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT53), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(KEYINPUT54), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT53), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n920), .B2(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n916), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n889), .A2(new_n890), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT115), .B(new_n788), .C1(new_n712), .C2(new_n714), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n896), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n929), .B1(new_n932), .B2(new_n899), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT54), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n927), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n925), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n878), .A2(new_n885), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(G952), .A2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n850), .B1(new_n937), .B2(new_n938), .ZN(G75));
  NAND2_X1  g753(.A1(new_n927), .A2(new_n933), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(G210), .A3(G902), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n379), .A2(new_n384), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n344), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT55), .Z(new_n944));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(KEYINPUT56), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n941), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n941), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n340), .A2(G952), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G51));
  NAND2_X1  g764(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n935), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n811), .B(KEYINPUT57), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n319), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n940), .A2(G902), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(new_n810), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n949), .B1(new_n955), .B2(new_n957), .ZN(G54));
  NAND2_X1  g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT122), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n524), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n949), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n940), .A2(G902), .A3(new_n520), .A4(new_n960), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(G60));
  INV_X1    g779(.A(new_n651), .ZN(new_n966));
  XNOR2_X1  g780(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n936), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n647), .A2(new_n649), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n968), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n925), .B2(new_n935), .ZN(new_n974));
  INV_X1    g788(.A(new_n971), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT124), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n971), .A2(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n949), .B1(new_n952), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(G63));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n895), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n900), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n801), .A2(new_n916), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n984), .A2(new_n926), .B1(new_n901), .B2(new_n929), .ZN(new_n985));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  OAI22_X1  g801(.A1(new_n985), .A2(new_n987), .B1(new_n623), .B2(new_n624), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n963), .ZN(new_n989));
  INV_X1    g803(.A(new_n685), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n985), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n980), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n991), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n993), .A2(new_n988), .A3(KEYINPUT61), .A4(new_n963), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n579), .B2(new_n342), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n922), .A2(new_n905), .A3(new_n902), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(G953), .ZN(new_n998));
  INV_X1    g812(.A(G898), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n942), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n998), .B(new_n1000), .Z(G69));
  NAND2_X1  g815(.A1(new_n427), .A2(new_n429), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(new_n516), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n930), .A2(new_n931), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n739), .A3(new_n744), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1006));
  OR3_X1    g820(.A1(new_n747), .A2(new_n790), .A3(new_n903), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n832), .B1(new_n718), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n839), .B2(new_n841), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT62), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1004), .A2(new_n739), .A3(new_n1010), .A4(new_n744), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1006), .A2(new_n1009), .A3(new_n340), .A4(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1003), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n286), .A2(G900), .A3(G953), .ZN(new_n1015));
  INV_X1    g829(.A(new_n801), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n913), .A2(new_n747), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n819), .A2(new_n710), .A3(new_n717), .A4(new_n1017), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n1016), .A2(new_n804), .A3(new_n832), .A4(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1004), .A2(new_n744), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1019), .A2(new_n842), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1014), .B1(new_n1022), .B2(new_n1003), .ZN(G72));
  NAND4_X1  g837(.A1(new_n1019), .A2(new_n1020), .A3(new_n842), .A4(new_n997), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  AND3_X1   g841(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1025), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n449), .A2(new_n436), .A3(new_n414), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n918), .A2(new_n924), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n464), .A2(KEYINPUT126), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n464), .A2(KEYINPUT126), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1033), .A2(new_n434), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n1027), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT127), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n949), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1006), .A2(new_n1009), .A3(new_n997), .A4(new_n1011), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1039), .A2(new_n1027), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n421), .B1(new_n430), .B2(new_n463), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1031), .A2(new_n1042), .ZN(G57));
endmodule


