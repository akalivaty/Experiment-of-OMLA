//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(new_n195), .B1(new_n192), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(KEYINPUT80), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n196), .B2(new_n197), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT81), .B(G101), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n200), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT2), .B(G113), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G119), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT67), .A3(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G119), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n211), .B1(new_n215), .B2(KEYINPUT69), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT68), .B(G116), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G119), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n205), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(KEYINPUT69), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n217), .A3(G119), .ZN(new_n222));
  INV_X1    g036(.A(new_n205), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n211), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(KEYINPUT70), .A3(new_n224), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n204), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n207), .A2(G119), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n221), .A2(new_n222), .A3(new_n211), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n232), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n224), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT82), .B1(new_n194), .B2(G104), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n192), .A3(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n194), .A2(G104), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT83), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n196), .A2(new_n202), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT83), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n245), .A3(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n190), .B1(new_n229), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n247), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n224), .A3(new_n235), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n220), .A2(KEYINPUT70), .A3(new_n224), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT70), .B1(new_n220), .B2(new_n224), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n251), .B(new_n189), .C1(new_n254), .C2(new_n204), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n255), .A3(KEYINPUT6), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT64), .A2(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT64), .A2(G146), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(KEYINPUT65), .B1(G143), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n260), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT64), .A2(G146), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(G143), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(G146), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(new_n257), .ZN(new_n276));
  OAI21_X1  g090(.A(G125), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n265), .A2(G143), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n268), .A3(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n262), .A2(new_n263), .A3(new_n261), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n286));
  OAI21_X1  g100(.A(G128), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n281), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G125), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G953), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G224), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n291), .B(new_n293), .Z(new_n294));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n295), .B(new_n190), .C1(new_n229), .C2(new_n248), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n256), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n189), .B(KEYINPUT8), .Z(new_n298));
  NAND2_X1  g112(.A1(new_n236), .A2(new_n247), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n251), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n277), .B2(new_n290), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n277), .A2(new_n290), .A3(new_n301), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n304), .B2(new_n255), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G210), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n297), .A2(new_n305), .A3(new_n307), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G140), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT79), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n292), .A2(G227), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n288), .A2(new_n247), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n278), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n280), .B1(new_n275), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n320), .A2(new_n244), .A3(new_n243), .A4(new_n246), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  INV_X1    g137(.A(G134), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G137), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT11), .A3(G134), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n327), .A3(new_n331), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT12), .B1(new_n333), .B2(KEYINPUT84), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n335), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n322), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n271), .B2(new_n272), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n283), .B1(new_n340), .B2(new_n267), .ZN(new_n341));
  INV_X1    g155(.A(new_n268), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n287), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n280), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n250), .A2(new_n344), .A3(KEYINPUT10), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n321), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n333), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n200), .A2(new_n201), .A3(new_n203), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n284), .A2(new_n259), .B1(new_n275), .B2(new_n257), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n347), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n317), .B1(new_n339), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n337), .B1(new_n322), .B2(new_n333), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n348), .B(new_n335), .C1(new_n318), .C2(new_n321), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n317), .B(new_n352), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n316), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n352), .A2(new_n315), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n333), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(G469), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n336), .A2(KEYINPUT86), .A3(new_n338), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n354), .B2(new_n355), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n366), .A3(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n352), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n316), .ZN(new_n369));
  AOI21_X1  g183(.A(G902), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G469), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(G469), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G221), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G902), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n261), .B2(G128), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n278), .A2(KEYINPUT89), .A3(G143), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n382), .A2(new_n383), .B1(G128), .B2(new_n261), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n384), .A2(new_n324), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT13), .B1(new_n382), .B2(new_n383), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT13), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n384), .B1(new_n388), .B2(new_n324), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT88), .B(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G116), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n218), .A2(G122), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n194), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n194), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n384), .B(new_n324), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n392), .A2(KEYINPUT14), .B1(G116), .B2(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n218), .A2(new_n400), .A3(G122), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n194), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n387), .A2(new_n396), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G217), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n376), .A2(new_n404), .A3(G953), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n399), .A2(new_n401), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n393), .B(new_n397), .C1(new_n408), .C2(new_n194), .ZN(new_n409));
  OAI221_X1 g223(.A(new_n389), .B1(new_n385), .B2(new_n386), .C1(new_n394), .C2(new_n395), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n289), .A2(KEYINPUT16), .A3(G140), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT78), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G125), .B(G140), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(G146), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G237), .A2(G953), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(G143), .A3(G214), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G143), .B1(new_n424), .B2(G214), .ZN(new_n427));
  OAI21_X1  g241(.A(G131), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n292), .A3(G214), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n261), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n331), .A3(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n262), .A2(new_n263), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n423), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n425), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT18), .A3(G131), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n420), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n265), .B2(new_n420), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT18), .A2(G131), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n431), .A2(new_n425), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(G113), .B(G122), .Z(new_n447));
  XOR2_X1   g261(.A(KEYINPUT87), .B(G104), .Z(new_n448));
  XOR2_X1   g262(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n449), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n439), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n433), .B2(KEYINPUT17), .ZN(new_n453));
  INV_X1    g267(.A(G140), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n289), .A2(G140), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT16), .ZN(new_n457));
  OR3_X1    g271(.A1(new_n289), .A2(KEYINPUT16), .A3(G140), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n422), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n265), .B1(new_n459), .B2(new_n418), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n423), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n451), .B(new_n445), .C1(new_n453), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n416), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT20), .B(new_n466), .C1(new_n450), .C2(new_n462), .ZN(new_n467));
  INV_X1    g281(.A(G475), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n445), .B1(new_n453), .B2(new_n461), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n449), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n465), .A2(new_n467), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n415), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n292), .A2(G952), .ZN(new_n475));
  INV_X1    g289(.A(G234), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n429), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT90), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n378), .B(new_n292), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n311), .A2(new_n374), .A3(new_n380), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n424), .A2(G210), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT26), .B(G101), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT73), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n326), .A2(G134), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n328), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n495), .B(G131), .C1(new_n494), .C2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n332), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n344), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n350), .A2(new_n333), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n227), .A2(new_n228), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n254), .A2(new_n499), .A3(new_n500), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT71), .B1(new_n288), .B2(new_n497), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT71), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n278), .B1(new_n273), .B2(KEYINPUT1), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n266), .B2(new_n268), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n498), .B(new_n508), .C1(new_n510), .C2(new_n281), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n500), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT72), .B1(new_n512), .B2(new_n502), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n497), .B1(new_n343), .B2(new_n280), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n514), .A2(new_n508), .B1(new_n333), .B2(new_n350), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n254), .A3(new_n516), .A4(new_n507), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n517), .A3(KEYINPUT28), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n492), .B1(new_n506), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n515), .B2(new_n507), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n499), .A2(new_n520), .A3(new_n500), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n502), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n513), .A2(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n491), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(new_n502), .B1(new_n513), .B2(new_n517), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT31), .A3(new_n491), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n519), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n487), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n519), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT31), .B1(new_n531), .B2(new_n491), .ZN(new_n538));
  AND4_X1   g352(.A1(KEYINPUT31), .A2(new_n524), .A3(new_n525), .A4(new_n491), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n531), .B2(new_n491), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n506), .A2(new_n518), .A3(new_n492), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n504), .A2(new_n505), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n513), .A2(new_n517), .B1(new_n502), .B2(new_n512), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(new_n505), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n491), .A2(KEYINPUT29), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n378), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G472), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n536), .A2(new_n541), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n209), .A2(G128), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n209), .A2(G128), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n553), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n556), .C1(new_n553), .C2(new_n563), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT77), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G110), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n461), .B(new_n560), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n557), .A2(new_n559), .B1(new_n566), .B2(G110), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n423), .A3(new_n441), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n375), .A2(new_n476), .A3(G953), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n576), .A3(new_n572), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n378), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n404), .B1(G234), .B2(new_n378), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n578), .A2(new_n579), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(G902), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n485), .A2(new_n552), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(new_n202), .Z(G3));
  OAI21_X1  g402(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n540), .A2(new_n534), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n374), .A2(new_n586), .A3(new_n380), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n297), .A2(new_n305), .A3(new_n307), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n307), .B1(new_n297), .B2(new_n305), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n187), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n403), .A2(new_n406), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT33), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n407), .A2(new_n600), .A3(new_n411), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(G478), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n413), .A2(new_n378), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n412), .B2(new_n413), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR4_X1   g419(.A1(new_n596), .A2(new_n473), .A3(new_n483), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n592), .A2(new_n593), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n610));
  INV_X1    g424(.A(new_n415), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n473), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n612), .B2(new_n483), .ZN(new_n613));
  INV_X1    g427(.A(new_n483), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n611), .A2(KEYINPUT91), .A3(new_n473), .A4(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n613), .A2(new_n311), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n592), .A3(new_n593), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NOR2_X1   g433(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n573), .B(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n582), .A2(new_n583), .B1(new_n585), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n485), .A2(new_n592), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT37), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  AND3_X1   g440(.A1(new_n536), .A2(new_n541), .A3(new_n551), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n477), .B(KEYINPUT92), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(G900), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n482), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n611), .A2(new_n473), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n622), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(new_n374), .A3(new_n311), .A4(new_n380), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT93), .B1(new_n627), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n374), .A2(new_n311), .A3(new_n380), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n552), .A3(new_n638), .A4(new_n634), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  AND2_X1   g455(.A1(new_n536), .A2(new_n541), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n547), .A2(new_n492), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n491), .B2(new_n531), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n644), .B2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n309), .A2(new_n310), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n611), .A2(new_n472), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n623), .A2(new_n188), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n631), .B(KEYINPUT39), .Z(new_n653));
  AND3_X1   g467(.A1(new_n374), .A2(new_n380), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT40), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT95), .B(G143), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G45));
  AND4_X1   g472(.A1(new_n472), .A2(new_n602), .A3(new_n604), .A4(new_n632), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n187), .C1(new_n594), .C2(new_n595), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT96), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n647), .A2(new_n662), .A3(new_n187), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n374), .A2(new_n380), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n552), .A3(new_n665), .A4(new_n623), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT97), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n374), .A2(new_n380), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n661), .B2(new_n663), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n552), .A4(new_n623), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n370), .B2(new_n371), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n370), .B2(KEYINPUT98), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n677), .B(G902), .C1(new_n367), .C2(new_n369), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n352), .A2(new_n315), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n354), .A2(new_n355), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(KEYINPUT86), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n682), .A2(new_n366), .B1(new_n316), .B2(new_n368), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n677), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n370), .A2(KEYINPUT98), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n674), .A4(G469), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n379), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n606), .A3(new_n552), .A4(new_n586), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n616), .A2(new_n687), .A3(new_n552), .A4(new_n586), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n311), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n552), .A2(new_n484), .A3(new_n623), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n209), .ZN(G21));
  AOI21_X1  g510(.A(new_n492), .B1(new_n548), .B2(KEYINPUT100), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n546), .C1(new_n547), .C2(new_n505), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n528), .A2(new_n532), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n535), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(G472), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n540), .B2(new_n378), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n647), .A2(new_n187), .A3(new_n614), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n650), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n687), .A3(new_n586), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  INV_X1    g523(.A(new_n659), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n702), .A2(new_n704), .A3(new_n622), .A4(new_n710), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n596), .B(new_n379), .C1(new_n679), .C2(new_n686), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NAND3_X1  g528(.A1(new_n309), .A2(new_n187), .A3(new_n310), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n668), .A2(new_n715), .A3(new_n716), .A4(new_n710), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT32), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n533), .B2(new_n535), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n541), .A3(new_n551), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n586), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n720), .B2(new_n586), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n717), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n668), .A2(new_n715), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n552), .A3(new_n586), .A4(new_n659), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n716), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  INV_X1    g543(.A(new_n633), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(new_n552), .A3(new_n586), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  INV_X1    g546(.A(new_n372), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n358), .A2(KEYINPUT45), .A3(new_n362), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT85), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n315), .B1(new_n737), .B2(new_n356), .ZN(new_n738));
  INV_X1    g552(.A(new_n362), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n734), .A2(new_n740), .A3(G469), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n373), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n733), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n373), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n380), .ZN(new_n747));
  INV_X1    g561(.A(new_n653), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT102), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n379), .B1(new_n744), .B2(new_n745), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n653), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n605), .B2(new_n472), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n473), .A2(new_n755), .A3(new_n602), .A4(new_n604), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT103), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n623), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n757), .B1(new_n754), .B2(new_n756), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n591), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  INV_X1    g577(.A(new_n715), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT44), .B1(new_n761), .B2(new_n591), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n753), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n747), .B2(KEYINPUT47), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n750), .A2(KEYINPUT105), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n747), .A2(new_n776), .A3(KEYINPUT47), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT106), .B1(new_n750), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n552), .A2(new_n715), .A3(new_n586), .A4(new_n710), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  AND2_X1   g596(.A1(new_n679), .A2(new_n686), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT49), .Z(new_n784));
  NAND3_X1  g598(.A1(new_n586), .A2(new_n187), .A3(new_n380), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n649), .A2(new_n472), .A3(new_n605), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n646), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n687), .A2(new_n764), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n756), .A2(new_n754), .A3(new_n629), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n722), .A2(new_n723), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n791), .B(new_n792), .C1(KEYINPUT115), .C2(KEYINPUT48), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(KEYINPUT115), .B2(KEYINPUT48), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n793), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n586), .A2(new_n787), .A3(new_n789), .A4(new_n478), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n605), .A2(new_n473), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n705), .A2(new_n586), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n790), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n798), .B(new_n475), .C1(new_n693), .C2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n794), .B(new_n795), .C1(new_n802), .C2(KEYINPUT114), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(KEYINPUT114), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n783), .A2(new_n380), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n775), .B2(new_n779), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n806), .A2(new_n715), .A3(new_n801), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n472), .B1(new_n602), .B2(new_n604), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n702), .A2(new_n704), .A3(new_n622), .ZN(new_n809));
  INV_X1    g623(.A(new_n791), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n796), .A2(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n687), .A2(new_n188), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT112), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n801), .A3(new_n649), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT50), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n817), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n807), .A2(new_n815), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n804), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n636), .A2(new_n639), .B1(new_n711), .B2(new_n712), .ZN(new_n825));
  INV_X1    g639(.A(new_n650), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n311), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n622), .A2(new_n632), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT110), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n646), .A2(new_n665), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n672), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n672), .A2(new_n825), .A3(KEYINPUT52), .A4(new_n831), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n728), .A2(new_n731), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n797), .A2(KEYINPUT107), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT107), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n605), .B2(new_n473), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n706), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n592), .A2(new_n842), .A3(new_n593), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n587), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT108), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT108), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n587), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n706), .A2(new_n612), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n592), .A2(new_n849), .A3(new_n593), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n708), .A2(new_n688), .A3(new_n624), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT109), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n700), .A2(new_n701), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n534), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n589), .A3(new_n623), .A4(new_n659), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n665), .A2(new_n764), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n809), .A2(new_n725), .A3(KEYINPUT109), .A4(new_n659), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n668), .A2(new_n474), .A3(new_n631), .A4(new_n715), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n627), .A2(new_n622), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n837), .A2(new_n848), .A3(new_n853), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n824), .B1(new_n836), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n853), .A2(new_n848), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n728), .A2(new_n863), .A3(new_n731), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n834), .A2(new_n835), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT53), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n868), .B2(new_n869), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n876), .A3(new_n870), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n823), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n788), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n292), .A2(G952), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n256), .A2(new_n296), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n294), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n871), .A2(G210), .A3(G902), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(G902), .B1(new_n873), .B2(new_n874), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n308), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n888), .B(KEYINPUT119), .Z(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n883), .B(new_n891), .C1(new_n895), .C2(new_n897), .ZN(G51));
  INV_X1    g712(.A(new_n741), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n899), .A3(new_n894), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n875), .A2(new_n877), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n373), .B(KEYINPUT57), .Z(new_n903));
  AOI21_X1  g717(.A(new_n683), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n900), .B2(KEYINPUT120), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n883), .B1(new_n901), .B2(new_n905), .ZN(G54));
  AND2_X1   g720(.A1(KEYINPUT58), .A2(G475), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n893), .A2(new_n894), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n462), .A3(new_n450), .ZN(new_n909));
  INV_X1    g723(.A(new_n883), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n893), .A2(new_n463), .A3(new_n894), .A4(new_n907), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G60));
  XNOR2_X1  g726(.A(new_n603), .B(KEYINPUT59), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n879), .A2(new_n872), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n599), .A2(new_n601), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n913), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n883), .B1(new_n902), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n873), .B2(new_n874), .ZN(new_n927));
  INV_X1    g741(.A(new_n584), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n883), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n871), .A2(new_n621), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  AOI21_X1  g753(.A(new_n292), .B1(new_n480), .B2(G224), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n866), .B2(new_n292), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n884), .B1(G898), .B2(new_n292), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(G69));
  AOI21_X1  g757(.A(new_n715), .B1(new_n841), .B2(new_n612), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n654), .A3(new_n552), .A4(new_n586), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n781), .A2(new_n769), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n656), .A2(new_n672), .A3(new_n825), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n656), .A2(new_n672), .A3(new_n825), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n292), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n530), .B(KEYINPUT124), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n435), .A2(new_n436), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n292), .B1(G227), .B2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n792), .A2(new_n827), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n753), .B1(new_n768), .B2(new_n959), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n672), .A2(new_n728), .A3(new_n731), .A4(new_n825), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n781), .A3(new_n961), .A4(new_n292), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n956), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n963), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n956), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n957), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n969), .B2(new_n957), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(KEYINPUT127), .B(new_n965), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OR2_X1    g793(.A1(new_n946), .A2(new_n951), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n866), .ZN(new_n981));
  INV_X1    g795(.A(new_n531), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n491), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n531), .B(new_n491), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n871), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n960), .A2(new_n781), .A3(new_n961), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n979), .B1(new_n986), .B2(new_n866), .ZN(new_n987));
  INV_X1    g801(.A(new_n491), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n988), .A3(new_n531), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n910), .A2(new_n983), .A3(new_n985), .A4(new_n989), .ZN(G57));
endmodule


