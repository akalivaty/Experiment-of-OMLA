//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT2), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  XNOR2_X1  g019(.A(G155gat), .B(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT74), .B(G155gat), .Z(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(KEYINPUT73), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(G141gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n221), .A4(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n223), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n215), .B1(new_n216), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G228gat), .ZN(new_n239));
  INV_X1    g038(.A(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n216), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n213), .B(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n237), .A2(KEYINPUT81), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n224), .B1(new_n237), .B2(KEYINPUT81), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n235), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n241), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(G22gat), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n241), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n223), .A2(new_n232), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n216), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT3), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n253), .B1(new_n234), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G22gat), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n246), .A2(new_n236), .A3(new_n241), .A4(new_n238), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n252), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n252), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n252), .A2(new_n262), .ZN(new_n267));
  INV_X1    g066(.A(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n202), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n262), .A3(new_n263), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT82), .B(G50gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n272), .A3(new_n274), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT27), .B(G183gat), .Z(new_n280));
  OAI21_X1  g079(.A(KEYINPUT67), .B1(new_n280), .B2(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT28), .A4(new_n285), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT26), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(new_n285), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT1), .ZN(new_n303));
  XOR2_X1   g102(.A(G127gat), .B(G134gat), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT64), .ZN(new_n307));
  NOR2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n293), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n293), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n285), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(new_n306), .C1(new_n311), .C2(KEYINPUT66), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n319), .B(new_n314), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n313), .A2(new_n318), .B1(new_n323), .B2(KEYINPUT25), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n305), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n305), .ZN(new_n326));
  INV_X1    g125(.A(new_n300), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n287), .B2(new_n291), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n318), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n326), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G227gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT34), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT34), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n325), .A2(new_n332), .A3(new_n337), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(new_n335), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n344), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n333), .B2(new_n335), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n336), .B(new_n338), .C1(new_n350), .C2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n348), .B1(new_n346), .B2(new_n351), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n279), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n346), .A2(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT86), .A3(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n236), .A2(new_n326), .A3(new_n233), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n305), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n223), .A2(new_n305), .A3(new_n232), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n365), .B2(new_n369), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n363), .B(new_n364), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n361), .A2(new_n369), .A3(new_n365), .A4(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n235), .A2(new_n326), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(new_n362), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n373), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT78), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n387), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n372), .B(new_n386), .C1(new_n378), .C2(new_n379), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G226gat), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n301), .B(new_n324), .C1(new_n398), .C2(new_n240), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n216), .B1(new_n398), .B2(new_n240), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n328), .B2(new_n331), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n245), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n401), .A3(new_n215), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT71), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n403), .A2(new_n412), .A3(new_n404), .A4(new_n408), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT35), .ZN(new_n415));
  INV_X1    g214(.A(new_n404), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n215), .B1(new_n399), .B2(new_n401), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n409), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n403), .A2(KEYINPUT30), .A3(new_n404), .A4(new_n408), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  AND4_X1   g220(.A1(new_n278), .A2(new_n360), .A3(new_n397), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n357), .A2(new_n352), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n276), .B2(new_n277), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n420), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n396), .B2(new_n388), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n415), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n376), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n375), .A2(new_n376), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(new_n431), .A3(new_n376), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n386), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT40), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n433), .A2(KEYINPUT40), .A3(new_n386), .A4(new_n434), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n393), .A3(new_n425), .A4(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n266), .A2(new_n272), .A3(new_n274), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n274), .B1(new_n266), .B2(new_n272), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n410), .A2(new_n413), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n404), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n403), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n404), .A2(new_n444), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT37), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n418), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n449), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n409), .B1(new_n405), .B2(KEYINPUT37), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n403), .B2(new_n404), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n443), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n392), .A2(new_n396), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n442), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n423), .B(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n278), .B2(new_n426), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n422), .A2(new_n427), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G1gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT16), .ZN(new_n466));
  INV_X1    g265(.A(G15gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G22gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n260), .A2(G15gat), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(G1gat), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g270(.A(G8gat), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n260), .A2(G15gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n467), .A2(G22gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G8gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(G43gat), .A2(G50gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(G43gat), .A2(G50gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT15), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n483), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G43gat), .ZN(new_n500));
  INV_X1    g299(.A(G50gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  NAND2_X1  g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n491), .A2(new_n484), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n483), .A3(new_n494), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n484), .A2(new_n485), .B1(new_n509), .B2(new_n490), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n493), .B1(new_n510), .B2(new_n487), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n483), .A3(new_n494), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n504), .A2(new_n503), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT89), .B(G43gat), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n511), .A2(new_n483), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n516), .A2(KEYINPUT90), .A3(new_n479), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT90), .B1(new_n516), .B2(new_n479), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT13), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n512), .A2(new_n515), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n470), .A2(new_n471), .A3(G8gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n523), .A2(new_n495), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(KEYINPUT90), .A3(new_n479), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n496), .B2(new_n507), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n523), .A2(new_n495), .A3(KEYINPUT17), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n480), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n520), .A2(KEYINPUT18), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(new_n534), .A3(new_n520), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n522), .A2(new_n537), .A3(KEYINPUT93), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(KEYINPUT92), .A3(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n540), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G169gat), .B(G197gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n544), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n522), .A2(new_n555), .A3(new_n537), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n464), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G71gat), .B(G78gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT20), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n573), .B(new_n574), .ZN(new_n580));
  INV_X1    g379(.A(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n579), .B2(new_n582), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n480), .B1(new_n571), .B2(new_n572), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n579), .A2(new_n582), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n583), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n590), .B1(new_n594), .B2(new_n585), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT95), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT41), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n602), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT97), .A2(G99gat), .A3(G106gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT97), .B1(G99gat), .B2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT8), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n601), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n601), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n602), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  OAI21_X1  g416(.A(G92gat), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n615), .B1(new_n618), .B2(new_n605), .ZN(new_n619));
  INV_X1    g418(.A(new_n610), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(KEYINPUT8), .A3(new_n608), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n613), .A2(KEYINPUT98), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(new_n601), .C1(new_n607), .C2(new_n612), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n600), .B1(new_n626), .B2(new_n516), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n625), .B(new_n623), .C1(new_n532), .C2(new_n533), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n598), .A2(new_n599), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT96), .Z(new_n635));
  XOR2_X1   g434(.A(G134gat), .B(G162gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n627), .A2(new_n628), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n630), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n642), .B2(new_n632), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n571), .A3(new_n625), .ZN(new_n645));
  INV_X1    g444(.A(new_n570), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n569), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n613), .A3(new_n622), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n649), .B(new_n653), .S(new_n654), .Z(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT102), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n654), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665));
  INV_X1    g464(.A(new_n654), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n649), .B2(new_n666), .ZN(new_n667));
  AOI211_X1 g466(.A(KEYINPUT101), .B(new_n654), .C1(new_n645), .C2(new_n648), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n667), .A2(new_n668), .A3(new_n658), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n660), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n596), .A2(new_n644), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n563), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n396), .A2(new_n388), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT103), .B(G1gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  AOI21_X1  g478(.A(new_n476), .B1(new_n674), .B2(new_n425), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n682));
  INV_X1    g481(.A(new_n563), .ZN(new_n683));
  INV_X1    g482(.A(new_n673), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n425), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT16), .B(G8gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n681), .A2(new_n682), .B1(KEYINPUT42), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(G1325gat));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n467), .A3(new_n360), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n563), .A2(new_n462), .A3(new_n673), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n467), .ZN(G1326gat));
  NOR3_X1   g496(.A1(new_n563), .A2(new_n278), .A3(new_n673), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n596), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n672), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n563), .A2(new_n644), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n489), .A3(new_n676), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(new_n644), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n464), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n464), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n522), .A2(KEYINPUT93), .A3(new_n537), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT93), .B1(new_n522), .B2(new_n537), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n541), .A2(KEYINPUT92), .A3(new_n543), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT92), .B1(new_n541), .B2(new_n543), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n555), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT107), .B1(new_n718), .B2(new_n560), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n557), .A2(new_n720), .A3(new_n561), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n702), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n711), .A2(new_n676), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n705), .B1(new_n489), .B2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n703), .A2(new_n490), .A3(new_n425), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT46), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n425), .A3(new_n723), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G36gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(G1329gat));
  INV_X1    g531(.A(new_n462), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n709), .A2(new_n733), .A3(new_n710), .A4(new_n723), .ZN(new_n734));
  INV_X1    g533(.A(new_n514), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n359), .A2(new_n735), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n703), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1330gat));
  NOR2_X1   g541(.A1(new_n440), .A2(new_n441), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n709), .A2(new_n743), .A3(new_n710), .A4(new_n723), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G50gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n703), .A2(new_n501), .A3(new_n743), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n701), .A2(new_n706), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n750), .A2(new_n671), .A3(new_n722), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n464), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n464), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n676), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n425), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT49), .B(G64gat), .Z(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n756), .B2(new_n462), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n360), .A2(new_n566), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n756), .A2(new_n278), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n567), .ZN(G1335gat));
  INV_X1    g569(.A(new_n722), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n596), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n671), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT112), .Z(new_n774));
  AND3_X1   g573(.A1(new_n711), .A2(new_n676), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n460), .A2(new_n463), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n355), .A2(new_n421), .A3(new_n358), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n277), .B2(new_n276), .ZN(new_n778));
  INV_X1    g577(.A(new_n423), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n426), .B(new_n779), .C1(new_n440), .C2(new_n441), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n778), .A2(new_n397), .B1(new_n780), .B2(KEYINPUT35), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n706), .B(new_n772), .C1(new_n776), .C2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n464), .A2(KEYINPUT51), .A3(new_n706), .A4(new_n772), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n676), .A2(new_n617), .A3(new_n671), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n775), .A2(new_n617), .B1(new_n786), .B2(new_n787), .ZN(G1336gat));
  NAND3_X1  g587(.A1(new_n784), .A2(KEYINPUT113), .A3(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n782), .A2(new_n790), .A3(new_n783), .ZN(new_n791));
  INV_X1    g590(.A(new_n425), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n792), .A2(G92gat), .A3(new_n672), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT114), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n789), .A2(new_n796), .A3(new_n791), .A4(new_n793), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n709), .A2(new_n425), .A3(new_n710), .A4(new_n774), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(new_n793), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n799), .B(new_n802), .C1(new_n786), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1337gat));
  NAND4_X1  g604(.A1(new_n709), .A2(new_n733), .A3(new_n710), .A4(new_n774), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  INV_X1    g606(.A(G99gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n360), .A2(new_n808), .A3(new_n671), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n786), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT115), .ZN(G1338gat));
  NAND4_X1  g610(.A1(new_n709), .A2(new_n743), .A3(new_n710), .A4(new_n774), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n278), .A2(G106gat), .A3(new_n672), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n813), .B(new_n814), .C1(new_n786), .C2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n789), .A2(new_n791), .A3(new_n815), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n814), .ZN(G1339gat));
  NAND3_X1  g619(.A1(new_n651), .A2(new_n652), .A3(new_n666), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n664), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n653), .A2(new_n825), .A3(new_n654), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n658), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n666), .B1(new_n653), .B2(new_n661), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n822), .B1(new_n830), .B2(new_n663), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n658), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n670), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n719), .A2(new_n721), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n519), .A2(new_n521), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n520), .B1(new_n530), .B2(new_n534), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n554), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n558), .B2(new_n559), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n670), .B2(new_n660), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n706), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n832), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n843), .A2(new_n824), .B1(new_n664), .B2(new_n669), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n831), .B2(new_n827), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n644), .A2(new_n839), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n644), .A2(new_n839), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n701), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n673), .B1(new_n719), .B2(new_n721), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n675), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n743), .A2(new_n425), .A3(new_n423), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n771), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n743), .B1(new_n854), .B2(new_n856), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n675), .A2(new_n425), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n360), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n562), .A2(G113gat), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  AOI21_X1  g667(.A(G120gat), .B1(new_n860), .B2(new_n671), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n360), .A2(G120gat), .A3(new_n671), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n864), .B2(new_n870), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n865), .B2(new_n701), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n701), .A2(G127gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n859), .B2(new_n873), .ZN(G1342gat));
  NOR3_X1   g673(.A1(new_n859), .A2(G134gat), .A3(new_n644), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n865), .B2(new_n644), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  AND2_X1   g677(.A1(new_n462), .A2(new_n863), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n840), .B1(new_n834), .B2(new_n562), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n849), .B(new_n852), .C1(new_n881), .C2(new_n706), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n855), .B1(new_n882), .B2(new_n701), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n276), .A2(KEYINPUT57), .A3(new_n277), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n850), .B1(new_n834), .B2(new_n851), .ZN(new_n887));
  AND4_X1   g686(.A1(new_n850), .A2(new_n851), .A3(new_n846), .A4(new_n844), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n560), .B1(new_n549), .B2(new_n556), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n841), .B1(new_n847), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n644), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n596), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT117), .B(new_n884), .C1(new_n893), .C2(new_n855), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n854), .A2(new_n856), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(new_n896), .B2(new_n743), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n879), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n792), .A2(new_n857), .A3(new_n743), .A4(new_n462), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n890), .A2(G141gat), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n904), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT118), .B(new_n879), .C1(new_n895), .C2(new_n897), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n771), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n906), .B1(new_n911), .B2(G141gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(new_n900), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n684), .A2(new_n890), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT121), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n891), .A2(new_n644), .B1(new_n834), .B2(new_n851), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n701), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n920), .B2(new_n743), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n885), .B1(new_n854), .B2(new_n856), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n879), .A2(new_n671), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n671), .A3(new_n909), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n230), .A2(KEYINPUT59), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n230), .A3(new_n671), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1345gat));
  NAND3_X1  g733(.A1(new_n901), .A2(new_n225), .A3(new_n596), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n910), .A2(new_n596), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n225), .ZN(G1346gat));
  AOI21_X1  g736(.A(G162gat), .B1(new_n901), .B2(new_n706), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n644), .A2(new_n226), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n910), .B2(new_n939), .ZN(G1347gat));
  AOI21_X1  g739(.A(new_n676), .B1(new_n854), .B2(new_n856), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(new_n425), .A3(new_n424), .ZN(new_n942));
  INV_X1    g741(.A(G169gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n771), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n676), .A2(new_n792), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(new_n359), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n862), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n890), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT123), .Z(G1348gat));
  INV_X1    g750(.A(G176gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n948), .A2(new_n952), .A3(new_n672), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n942), .A2(new_n671), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n952), .ZN(G1349gat));
  INV_X1    g754(.A(new_n948), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n298), .B1(new_n956), .B2(new_n596), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n596), .A2(new_n289), .A3(new_n290), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n942), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n956), .A2(new_n706), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(G190gat), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n961), .A3(G190gat), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n964), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n942), .A2(new_n285), .A3(new_n706), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1351gat));
  NAND4_X1  g772(.A1(new_n941), .A2(new_n425), .A3(new_n743), .A4(new_n462), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n771), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n923), .A2(new_n733), .A3(new_n946), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n562), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n671), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  AOI21_X1  g780(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n975), .A2(new_n671), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n975), .A2(new_n205), .A3(new_n596), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n946), .A2(new_n733), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n596), .B(new_n988), .C1(new_n921), .C2(new_n922), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n206), .A3(new_n706), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n706), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n993), .B1(new_n995), .B2(new_n206), .ZN(G1355gat));
endmodule


