//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT78), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n203), .A2(new_n204), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n205), .A2(new_n207), .A3(G146), .ZN(new_n224));
  INV_X1    g038(.A(new_n198), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n224), .A2(G128), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT80), .ZN(new_n229));
  INV_X1    g043(.A(new_n223), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G143), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n198), .B1(new_n231), .B2(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n231), .B2(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(G128), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n227), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n211), .A2(new_n237), .A3(new_n223), .A4(new_n227), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n244), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n239), .A2(KEYINPUT12), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n250), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT12), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n239), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n250), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n217), .A2(new_n220), .A3(new_n213), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G101), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n263), .A3(G101), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n205), .A2(new_n207), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n209), .ZN(new_n271));
  INV_X1    g085(.A(new_n210), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n224), .A2(new_n225), .A3(new_n267), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n259), .A2(new_n236), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n208), .A2(new_n210), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n200), .A2(new_n202), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n204), .B1(new_n278), .B2(new_n225), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n227), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n230), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT79), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n259), .B1(new_n211), .B2(new_n227), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n230), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n250), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n196), .B1(new_n258), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n196), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n276), .A2(new_n286), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n291), .B2(KEYINPUT82), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n276), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n190), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G469), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n281), .A2(KEYINPUT79), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n284), .B1(new_n283), .B2(new_n230), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n236), .A2(new_n259), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n265), .A2(new_n275), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT82), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n250), .A3(new_n294), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n288), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n195), .ZN(new_n307));
  INV_X1    g121(.A(new_n290), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n258), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G469), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n297), .A2(KEYINPUT83), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n313), .A3(G469), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n189), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n204), .A2(G119), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT24), .B(G110), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT71), .B1(new_n204), .B2(G119), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT72), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n318), .A3(new_n319), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n321), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT16), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n329), .A3(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n209), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(G146), .A3(new_n335), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n319), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n317), .A2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G110), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n326), .A2(new_n321), .ZN(new_n348));
  INV_X1    g162(.A(G110), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n341), .A2(new_n343), .A3(new_n349), .A4(new_n342), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n333), .A2(KEYINPUT73), .A3(G146), .A4(new_n335), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n330), .A2(new_n332), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n209), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n351), .A2(new_n353), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n346), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n347), .B1(new_n346), .B2(new_n357), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT74), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n346), .A2(new_n347), .A3(new_n357), .A4(new_n363), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n190), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(new_n190), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n324), .A2(new_n327), .ZN(new_n373));
  INV_X1    g187(.A(new_n338), .ZN(new_n374));
  AOI21_X1  g188(.A(G146), .B1(new_n333), .B2(new_n335), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n345), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n357), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n346), .A2(new_n347), .A3(new_n357), .ZN(new_n379));
  INV_X1    g193(.A(new_n363), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n381), .B2(new_n365), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT76), .B1(new_n382), .B2(KEYINPUT25), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n369), .B(G902), .C1(new_n381), .C2(new_n365), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n370), .B(new_n372), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n365), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n372), .A2(G902), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n232), .A2(new_n267), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n267), .A2(new_n268), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n208), .B2(new_n210), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n250), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G113), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n394), .A2(KEYINPUT2), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(KEYINPUT2), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n317), .A2(G116), .ZN(new_n398));
  INV_X1    g212(.A(G116), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G119), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n398), .B(new_n400), .C1(new_n395), .C2(new_n396), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n271), .A2(new_n272), .ZN(new_n406));
  OAI21_X1  g220(.A(G128), .B1(new_n226), .B2(new_n198), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n278), .A2(new_n204), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n406), .A2(new_n407), .B1(new_n232), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT65), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n241), .B2(G137), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n243), .A2(KEYINPUT65), .A3(G134), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n245), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G131), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n249), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n393), .B(new_n405), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT28), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n414), .A2(new_n249), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n280), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n405), .A4(new_n393), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT67), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n409), .B2(new_n415), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n280), .A2(new_n418), .A3(KEYINPUT67), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n393), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n417), .A2(new_n421), .B1(new_n425), .B2(new_n404), .ZN(new_n426));
  INV_X1    g240(.A(G237), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n191), .A3(G210), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT27), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G101), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT68), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n417), .A2(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n393), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT67), .B1(new_n280), .B2(new_n418), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n404), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n438));
  INV_X1    g252(.A(new_n431), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n434), .B2(new_n435), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n404), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n416), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n439), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n444), .A2(KEYINPUT31), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT31), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n432), .B(new_n440), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(G472), .A2(G902), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(KEYINPUT32), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT70), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n437), .B2(new_n439), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n431), .B1(new_n444), .B2(new_n416), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n419), .A2(new_n393), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n404), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n417), .B2(new_n421), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n439), .A2(new_n456), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n190), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT29), .B1(new_n426), .B2(new_n431), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n425), .B2(new_n441), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n445), .B1(new_n470), .B2(new_n404), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n468), .B(KEYINPUT70), .C1(new_n431), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G472), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n389), .B1(new_n454), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n187), .A2(new_n371), .A3(G953), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n399), .A2(G122), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n219), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n197), .B2(G128), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n204), .A2(KEYINPUT88), .A3(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(new_n486), .A3(new_n241), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n241), .B1(new_n485), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n478), .B2(G116), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT89), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n492), .A3(KEYINPUT14), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n399), .A2(G122), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT14), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n478), .A2(G116), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n219), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G107), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n481), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n485), .A2(new_n486), .A3(new_n241), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n486), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n231), .A2(KEYINPUT13), .A3(G128), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n485), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(G134), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n477), .B1(new_n500), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n494), .A2(new_n498), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G107), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n481), .C1(new_n487), .C2(new_n488), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(G134), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n503), .A3(new_n502), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n515), .A3(new_n476), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT90), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n513), .A2(new_n515), .A3(new_n518), .A4(new_n476), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n190), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT91), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n517), .A2(new_n519), .A3(new_n522), .A4(new_n190), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G478), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n520), .B2(KEYINPUT91), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n355), .B(KEYINPUT19), .Z(new_n532));
  NAND3_X1  g346(.A1(new_n427), .A2(new_n191), .A3(G214), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n231), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n427), .A2(new_n191), .A3(G143), .A4(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n248), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n532), .A2(G146), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n353), .A2(new_n354), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n355), .B(new_n209), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n534), .B(new_n535), .C1(new_n543), .C2(new_n248), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(G131), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n543), .ZN(new_n546));
  XNOR2_X1  g360(.A(G113), .B(G122), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(new_n212), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n537), .A2(KEYINPUT17), .A3(new_n538), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n337), .B(new_n338), .C1(new_n545), .C2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n546), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n541), .A2(new_n550), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NOR2_X1   g370(.A1(G475), .A2(G902), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n548), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n549), .B(new_n546), .C1(new_n539), .C2(new_n540), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT20), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n564), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n190), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n558), .A2(new_n562), .B1(new_n567), .B2(G475), .ZN(new_n568));
  INV_X1    g382(.A(new_n526), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n521), .B2(new_n523), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT92), .B1(new_n570), .B2(new_n529), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n531), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G214), .B1(G237), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G210), .B1(G237), .B2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT85), .B(G224), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT7), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n331), .B(new_n227), .C1(new_n277), .C2(new_n279), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n331), .B1(new_n390), .B2(new_n392), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT5), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G113), .B1(new_n398), .B2(KEYINPUT5), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n403), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n223), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n585), .B(G113), .C1(KEYINPUT5), .C2(new_n398), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(new_n216), .A3(new_n222), .A4(new_n403), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT8), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G125), .B1(new_n273), .B2(new_n274), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n596), .A2(KEYINPUT7), .A3(new_n579), .A4(new_n581), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n584), .A2(new_n595), .A3(new_n597), .A4(KEYINPUT86), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n262), .A2(new_n264), .A3(new_n404), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n593), .A3(new_n591), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n581), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(new_n580), .B1(new_n592), .B2(new_n594), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT86), .B1(new_n603), .B2(new_n597), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n190), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n591), .ZN(new_n606));
  INV_X1    g420(.A(new_n593), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT84), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT6), .A4(new_n600), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n602), .B(new_n578), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(KEYINPUT6), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n576), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n584), .A2(new_n595), .A3(new_n597), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n600), .A3(new_n598), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n190), .A3(new_n620), .A4(new_n575), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n574), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G952), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(G953), .ZN(new_n624));
  INV_X1    g438(.A(G234), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n427), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n190), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT21), .B(G898), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n572), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n315), .A2(new_n475), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  INV_X1    g449(.A(new_n388), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n367), .A2(new_n369), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n382), .A2(KEYINPUT25), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(KEYINPUT76), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n372), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT25), .B1(new_n386), .B2(new_n190), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n368), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n636), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n450), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n444), .A2(new_n446), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT31), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n444), .A2(KEYINPUT31), .A3(new_n446), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT68), .B(new_n431), .C1(new_n433), .C2(new_n436), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n644), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n449), .A2(new_n190), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(G472), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n315), .A2(new_n643), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n657));
  NAND3_X1  g471(.A1(new_n517), .A2(new_n519), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT94), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT94), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n517), .A2(new_n519), .A3(new_n660), .A4(new_n657), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT95), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n516), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n510), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n662), .B(new_n477), .C1(new_n500), .C2(new_n509), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(KEYINPUT33), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n525), .A2(G902), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n659), .A2(new_n661), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT96), .B(G478), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n520), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n558), .A2(new_n562), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n567), .A2(G475), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT97), .B1(new_n632), .B2(new_n675), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n574), .B(new_n630), .C1(new_n615), .C2(new_n621), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n674), .A4(new_n671), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n656), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  AOI21_X1  g499(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n570), .A2(KEYINPUT92), .A3(new_n529), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n677), .B(new_n568), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n656), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT35), .B(G107), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  XOR2_X1   g505(.A(new_n377), .B(KEYINPUT99), .Z(new_n692));
  NOR2_X1   g506(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n639), .A2(new_n642), .B1(new_n694), .B2(new_n387), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n615), .A2(new_n621), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n573), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n531), .A2(new_n571), .A3(new_n568), .A4(new_n631), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n315), .A2(new_n655), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  NAND2_X1  g517(.A1(new_n694), .A2(new_n387), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n385), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n622), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n454), .B2(new_n474), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n628), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n626), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n568), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n531), .B2(new_n571), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n315), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  XNOR2_X1  g528(.A(new_n710), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n315), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT40), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n674), .A2(new_n573), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n531), .B2(new_n571), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n695), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT100), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n447), .A2(new_n448), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n432), .A2(new_n440), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT32), .B(new_n450), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n471), .A2(new_n439), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n416), .A2(new_n439), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n190), .B1(new_n462), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n724), .B(new_n728), .C1(new_n653), .C2(new_n452), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n696), .B(KEYINPUT38), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n717), .A2(new_n721), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n231), .B(KEYINPUT101), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G45));
  NAND3_X1  g549(.A1(new_n671), .A2(new_n674), .A3(new_n710), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n315), .A2(new_n707), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  AOI21_X1  g553(.A(new_n196), .B1(new_n305), .B2(new_n288), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT12), .B1(new_n239), .B2(new_n250), .ZN(new_n741));
  INV_X1    g555(.A(new_n251), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(KEYINPUT81), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n290), .B1(new_n743), .B2(new_n253), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n190), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G469), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n311), .B(new_n190), .C1(new_n740), .C2(new_n744), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n188), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n475), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n681), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT41), .B(G113), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n688), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n399), .ZN(G18));
  OAI21_X1  g570(.A(new_n724), .B1(new_n653), .B2(new_n452), .ZN(new_n757));
  INV_X1    g571(.A(G472), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n468), .B1(new_n431), .B2(new_n471), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n466), .B1(new_n759), .B2(new_n455), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n760), .B2(new_n472), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n705), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n748), .A2(new_n749), .A3(new_n697), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n700), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G119), .ZN(G21));
  AOI211_X1 g580(.A(KEYINPUT104), .B(new_n636), .C1(new_n639), .C2(new_n642), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n385), .B2(new_n388), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n463), .A2(new_n431), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n647), .B2(new_n648), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT102), .B1(new_n772), .B2(new_n644), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT102), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(new_n450), .C1(new_n722), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT103), .B(G472), .Z(new_n777));
  NAND2_X1  g591(.A1(new_n654), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n770), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n746), .A2(new_n188), .A3(new_n747), .A4(new_n631), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n568), .A2(new_n574), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n696), .C1(new_n686), .C2(new_n687), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G122), .ZN(G24));
  NOR4_X1   g600(.A1(new_n748), .A2(new_n749), .A3(new_n697), .A4(new_n736), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n773), .A2(new_n775), .B1(new_n654), .B2(new_n777), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(KEYINPUT105), .A3(new_n705), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT105), .B1(new_n788), .B2(new_n705), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  INV_X1    g606(.A(KEYINPUT106), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n653), .B2(KEYINPUT32), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n449), .A2(new_n450), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT32), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(KEYINPUT106), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n724), .A3(new_n797), .A4(new_n474), .ZN(new_n798));
  INV_X1    g612(.A(new_n769), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n643), .A2(new_n768), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n749), .B1(new_n297), .B2(new_n747), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n615), .A2(new_n621), .A3(new_n573), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n736), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n806), .B(new_n643), .C1(new_n757), .C2(new_n761), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n802), .A2(new_n804), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n805), .A2(KEYINPUT42), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G131), .ZN(G33));
  INV_X1    g625(.A(new_n803), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n475), .A2(new_n712), .A3(new_n802), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  AOI21_X1  g628(.A(new_n674), .B1(new_n670), .B2(new_n668), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT43), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n817), .A2(new_n655), .A3(new_n695), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n803), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n204), .B1(new_n271), .B2(KEYINPUT1), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n227), .B1(new_n822), .B2(new_n232), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n823), .A2(new_n230), .B1(new_n228), .B2(KEYINPUT80), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n287), .B1(new_n824), .B2(new_n238), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n257), .B1(new_n825), .B2(KEYINPUT12), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT81), .B1(new_n825), .B2(KEYINPUT12), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n288), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n195), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n305), .A2(new_n308), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(KEYINPUT45), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT45), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n289), .B2(new_n295), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n833), .A3(G469), .ZN(new_n834));
  NAND2_X1  g648(.A1(G469), .A2(G902), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT46), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n311), .B2(new_n310), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(KEYINPUT46), .A3(new_n835), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n749), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n715), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n821), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT108), .B(G137), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G39));
  XNOR2_X1  g657(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n452), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n795), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n474), .A2(new_n849), .A3(new_n724), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n643), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n804), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(G140), .ZN(G42));
  NOR2_X1   g667(.A1(new_n817), .A2(new_n626), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n780), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n574), .A3(new_n732), .A4(new_n750), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n189), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n748), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n812), .B(new_n855), .C1(new_n847), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n748), .A2(new_n749), .A3(new_n803), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n776), .A2(new_n705), .A3(new_n778), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT105), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n788), .A2(KEYINPUT105), .A3(new_n705), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n864), .A2(new_n643), .A3(new_n627), .A4(new_n730), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n674), .A3(new_n671), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT51), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n798), .A2(new_n801), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  OAI21_X1  g691(.A(new_n624), .B1(new_n871), .B2(new_n675), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n855), .B2(new_n764), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT112), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n881), .B2(new_n873), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n877), .B(new_n879), .C1(new_n883), .C2(new_n862), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n720), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n696), .A2(new_n710), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n729), .A3(new_n802), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n791), .A2(new_n713), .A3(new_n738), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n868), .A2(new_n869), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n850), .A2(new_n698), .A3(new_n712), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n892), .A2(new_n787), .B1(new_n893), .B2(new_n315), .ZN(new_n894));
  AOI21_X1  g708(.A(G902), .B1(new_n829), .B2(new_n830), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT83), .B1(new_n895), .B2(new_n311), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n314), .A3(new_n747), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n859), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n698), .B(new_n737), .C1(new_n757), .C2(new_n761), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n729), .A2(new_n719), .A3(new_n695), .A4(new_n887), .ZN(new_n900));
  INV_X1    g714(.A(new_n802), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n898), .A2(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n891), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT111), .B1(new_n890), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n892), .A2(new_n809), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n527), .A2(new_n530), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n803), .A3(new_n711), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n763), .A2(new_n315), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n810), .A2(new_n813), .A3(new_n906), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n762), .A2(new_n699), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n911), .A2(new_n764), .B1(new_n780), .B2(new_n784), .ZN(new_n912));
  INV_X1    g726(.A(new_n688), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n475), .B(new_n750), .C1(new_n680), .C2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n634), .A3(new_n701), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT110), .B1(new_n671), .B2(new_n674), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT110), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n675), .A2(new_n917), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n916), .B(new_n918), .C1(new_n568), .C2(new_n907), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n656), .A2(new_n919), .A3(new_n632), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n910), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT111), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n894), .A2(new_n903), .A3(new_n891), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n905), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n921), .A2(KEYINPUT53), .A3(new_n924), .A4(new_n922), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n805), .A2(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n808), .A2(new_n809), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n813), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n906), .A2(new_n909), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n914), .A2(new_n765), .A3(new_n634), .A4(new_n785), .ZN(new_n937));
  INV_X1    g751(.A(new_n701), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n920), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n922), .A2(new_n924), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n927), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n926), .B2(new_n927), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n931), .B1(KEYINPUT54), .B2(new_n944), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n885), .A2(new_n945), .B1(new_n623), .B2(new_n191), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n748), .B(KEYINPUT49), .Z(new_n948));
  NAND4_X1  g762(.A1(new_n732), .A2(new_n859), .A3(new_n573), .A4(new_n815), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n948), .A2(new_n950), .A3(new_n730), .A4(new_n801), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT113), .ZN(new_n953));
  INV_X1    g767(.A(new_n951), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(G75));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n928), .A2(new_n930), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(G902), .ZN(new_n959));
  INV_X1    g773(.A(G210), .ZN(new_n960));
  OAI211_X1 g774(.A(KEYINPUT114), .B(new_n957), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n610), .A2(new_n613), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(new_n611), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n191), .A2(G952), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n961), .A2(new_n964), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT115), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n965), .A2(KEYINPUT115), .A3(new_n967), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(G51));
  INV_X1    g787(.A(KEYINPUT118), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT117), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n959), .B2(new_n834), .ZN(new_n976));
  INV_X1    g790(.A(new_n834), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n958), .A2(KEYINPUT117), .A3(G902), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n740), .A2(new_n744), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n835), .B(KEYINPUT57), .Z(new_n981));
  AOI21_X1  g795(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n931), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n983), .B2(KEYINPUT116), .ZN(new_n984));
  INV_X1    g798(.A(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n941), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT53), .B1(new_n987), .B2(new_n925), .ZN(new_n988));
  INV_X1    g802(.A(new_n930), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT54), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT116), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n979), .B1(new_n984), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n974), .B1(new_n995), .B2(new_n966), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n976), .A2(new_n978), .ZN(new_n997));
  INV_X1    g811(.A(new_n980), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n992), .B2(new_n993), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(KEYINPUT118), .A3(new_n967), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n996), .A2(new_n1002), .ZN(G54));
  INV_X1    g817(.A(new_n959), .ZN(new_n1004));
  AND2_X1   g818(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n555), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT119), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n966), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT119), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1004), .A2(new_n1010), .A3(new_n555), .A4(new_n1005), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT120), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT120), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1008), .A2(new_n1009), .A3(new_n1014), .A4(new_n1011), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G60));
  NAND3_X1  g830(.A1(new_n659), .A2(new_n661), .A3(new_n666), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G478), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT59), .Z(new_n1019));
  AOI211_X1 g833(.A(new_n1017), .B(new_n1019), .C1(new_n990), .C2(new_n991), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT121), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n945), .B2(new_n1019), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1021), .A2(new_n967), .A3(new_n1022), .ZN(G63));
  NOR2_X1   g837(.A1(new_n988), .A2(new_n989), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT60), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n967), .B1(new_n1027), .B2(new_n386), .ZN(new_n1028));
  INV_X1    g842(.A(new_n694), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1024), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT61), .ZN(new_n1031));
  OAI22_X1  g845(.A1(new_n1028), .A2(new_n1030), .B1(KEYINPUT122), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(KEYINPUT122), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1032), .B(new_n1033), .ZN(G66));
  OAI21_X1  g848(.A(G953), .B1(new_n577), .B2(new_n629), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n915), .A2(new_n920), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(G953), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n962), .B1(G898), .B2(new_n191), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G69));
  AOI21_X1  g853(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT124), .ZN(new_n1041));
  OR3_X1    g855(.A1(new_n840), .A2(new_n783), .A3(new_n875), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n852), .A2(new_n810), .A3(new_n813), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n894), .A2(new_n738), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n841), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n841), .A2(KEYINPUT126), .A3(new_n1045), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n191), .B(new_n1044), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n470), .B(new_n532), .Z(new_n1051));
  NAND2_X1  g865(.A1(G900), .A2(G953), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1053), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n733), .A2(new_n1045), .ZN(new_n1055));
  OR2_X1    g869(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n475), .A2(new_n812), .ZN(new_n1058));
  NOR3_X1   g872(.A1(new_n716), .A2(new_n919), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n841), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n1056), .A2(new_n852), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1051), .B1(new_n1061), .B2(new_n191), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n1041), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1041), .B(KEYINPUT125), .Z(new_n1064));
  INV_X1    g878(.A(KEYINPUT123), .ZN(new_n1065));
  OAI211_X1 g879(.A(new_n1053), .B(new_n1064), .C1(new_n1062), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g880(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(G72));
  NAND2_X1  g882(.A1(G472), .A2(G902), .ZN(new_n1069));
  XOR2_X1   g883(.A(new_n1069), .B(KEYINPUT63), .Z(new_n1070));
  INV_X1    g884(.A(new_n1036), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1070), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1072), .A2(new_n725), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n645), .B1(new_n471), .B2(new_n431), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n944), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g890(.A(new_n1036), .B(new_n1044), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1077));
  AND2_X1   g891(.A1(new_n1077), .A2(new_n1070), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n444), .A2(new_n416), .A3(new_n439), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n967), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g894(.A(KEYINPUT127), .ZN(new_n1081));
  NAND2_X1  g895(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g896(.A(KEYINPUT127), .B(new_n967), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n1076), .B1(new_n1082), .B2(new_n1083), .ZN(G57));
endmodule


