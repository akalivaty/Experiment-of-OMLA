//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1336, new_n1337, new_n1338, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  AND2_X1   g0023(.A1(KEYINPUT65), .A2(G77), .ZN(new_n224));
  NOR2_X1   g0024(.A1(KEYINPUT65), .A2(G77), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT66), .B(G244), .Z(new_n227));
  OAI211_X1 g0027(.A(new_n222), .B(new_n223), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT67), .Z(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT80), .ZN(new_n249));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  OR3_X1    g0052(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n250), .A2(new_n207), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n215), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G68), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n206), .B2(G20), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n253), .A2(new_n254), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT68), .B1(new_n262), .B2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(new_n207), .A3(G33), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n202), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n207), .A2(new_n262), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n268), .A2(new_n219), .B1(new_n207), .B2(G68), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n257), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT11), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n261), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  INV_X1    g0076(.A(G232), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G226), .B2(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G97), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n279), .A2(new_n283), .B1(new_n262), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n285), .A2(new_n286), .B1(G238), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AND2_X1   g0093(.A1(G1), .A2(G13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(KEYINPUT73), .A3(new_n289), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n291), .A2(new_n292), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n292), .B1(new_n291), .B2(new_n301), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n276), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n299), .A2(new_n300), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G226), .A2(G1698), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n277), .B2(G1698), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT3), .B(G33), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(G33), .B2(G97), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n294), .A2(new_n295), .ZN(new_n310));
  INV_X1    g0110(.A(G238), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT13), .B1(new_n305), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n291), .A2(new_n292), .A3(new_n301), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G179), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n292), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n305), .B2(new_n314), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n316), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n276), .B1(new_n321), .B2(G169), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n275), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(G200), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n315), .A2(G190), .A3(new_n316), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n274), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT75), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n219), .B1(new_n206), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n258), .A2(new_n328), .B1(new_n219), .B2(new_n255), .ZN(new_n329));
  INV_X1    g0129(.A(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT8), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT8), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G58), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n263), .A2(new_n265), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G150), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n201), .A2(new_n207), .B1(new_n268), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n257), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT72), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT72), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n341), .B(KEYINPUT9), .C1(new_n329), .C2(new_n337), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G222), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G223), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n308), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n283), .A2(new_n226), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n286), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n297), .B1(new_n313), .B2(new_n220), .ZN(new_n351));
  OAI21_X1  g0151(.A(G200), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n351), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G190), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT9), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT10), .B1(new_n343), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n329), .A2(new_n337), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n341), .B1(new_n358), .B2(KEYINPUT9), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n339), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n352), .A2(new_n355), .A3(new_n354), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n350), .A2(new_n351), .A3(G179), .ZN(new_n366));
  AOI21_X1  g0166(.A(G169), .B1(new_n353), .B2(new_n349), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n366), .A2(new_n367), .A3(new_n358), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT69), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n277), .A2(G1698), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n308), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n308), .B2(new_n372), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n308), .A2(G238), .A3(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n283), .A2(G107), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n286), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n297), .B1(new_n313), .B2(new_n227), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n370), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n257), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n266), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n224), .A2(new_n225), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n331), .A2(new_n333), .ZN(new_n388));
  INV_X1    g0188(.A(new_n268), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n387), .A2(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n384), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT70), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n387), .B2(new_n252), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n226), .A2(new_n255), .A3(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n258), .B(G77), .C1(G1), .C2(new_n207), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT71), .B1(new_n383), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n391), .A2(new_n397), .ZN(new_n401));
  INV_X1    g0201(.A(new_n379), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n308), .A2(new_n372), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT69), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n373), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n381), .B1(new_n406), .B2(new_n286), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n400), .B(new_n401), .C1(new_n407), .C2(new_n370), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(G190), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n380), .A2(new_n382), .ZN(new_n411));
  INV_X1    g0211(.A(G169), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G179), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n415), .A3(new_n398), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n365), .A2(new_n369), .A3(new_n410), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n388), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n206), .B2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n258), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n252), .B2(new_n388), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n330), .A2(new_n259), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n389), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(G20), .B1(new_n280), .B2(new_n282), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(KEYINPUT7), .B1(new_n308), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(G68), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n384), .B1(new_n430), .B2(KEYINPUT16), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n281), .B2(G33), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n262), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n282), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT7), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n308), .B2(G20), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n259), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n432), .B1(new_n440), .B2(new_n426), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n421), .B1(new_n431), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n310), .A2(G232), .A3(new_n312), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n297), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G87), .ZN(new_n445));
  OR2_X1    g0245(.A1(G223), .A2(G1698), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n220), .A2(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n448), .B2(new_n283), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n286), .ZN(new_n450));
  INV_X1    g0250(.A(G190), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n444), .A2(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n370), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n444), .A2(new_n450), .A3(new_n456), .A4(new_n451), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n442), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n454), .A2(G169), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n444), .A2(new_n450), .A3(G179), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n442), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n442), .A2(new_n458), .A3(KEYINPUT17), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n419), .A2(new_n258), .B1(new_n255), .B2(new_n418), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n424), .A2(new_n425), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n428), .B1(new_n280), .B2(new_n282), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n283), .A2(new_n207), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(new_n438), .ZN(new_n472));
  OAI211_X1 g0272(.A(KEYINPUT16), .B(new_n469), .C1(new_n472), .C2(new_n259), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n257), .ZN(new_n474));
  INV_X1    g0274(.A(new_n432), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT77), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n428), .B1(new_n478), .B2(new_n435), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n480));
  OAI21_X1  g0280(.A(G68), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n475), .B1(new_n481), .B2(new_n469), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n468), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n463), .B1(new_n414), .B2(new_n454), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n462), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n461), .A2(new_n466), .A3(new_n467), .A4(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n327), .A2(new_n417), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n323), .A2(KEYINPUT75), .A3(new_n326), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n249), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n416), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n401), .B1(new_n407), .B2(new_n370), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(KEYINPUT71), .B1(G190), .B2(new_n407), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n408), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n466), .A2(new_n487), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT17), .B1(new_n442), .B2(new_n458), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n368), .B1(new_n357), .B2(new_n364), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n497), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NOR4_X1   g0302(.A1(new_n502), .A2(new_n490), .A3(new_n327), .A4(KEYINPUT80), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT82), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n206), .A2(G45), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G41), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT82), .A3(new_n206), .A4(G45), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(G41), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(G257), .A3(new_n310), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n206), .B(G45), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n516), .B2(new_n505), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n296), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(new_n345), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT4), .A2(G244), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(G1698), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n308), .A2(new_n525), .B1(G33), .B2(G283), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n310), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n370), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n286), .B1(new_n517), .B2(new_n511), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n530));
  AOI22_X1  g0330(.A1(G257), .A2(new_n529), .B1(new_n530), .B2(new_n296), .ZN(new_n531));
  INV_X1    g0331(.A(new_n527), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n528), .B1(new_n533), .B2(G190), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n479), .B2(new_n480), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n537), .A2(new_n284), .A3(G107), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G20), .B1(G77), .B2(new_n389), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n384), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n252), .A2(G97), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n257), .B(new_n255), .C1(new_n206), .C2(G33), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT81), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n437), .B2(new_n439), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n539), .B1(new_n537), .B2(new_n536), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n551), .A2(new_n207), .B1(new_n202), .B2(new_n268), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n257), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT81), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n546), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n534), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n532), .A2(new_n414), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT83), .B1(new_n557), .B2(new_n519), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n546), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n531), .A2(new_n560), .A3(new_n414), .A4(new_n532), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n412), .B1(new_n519), .B2(new_n527), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT84), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n308), .A2(new_n207), .A3(G68), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n284), .B1(new_n263), .B2(new_n265), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(KEYINPUT19), .ZN(new_n570));
  NAND3_X1  g0370(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n571), .A2(KEYINPUT86), .A3(new_n207), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT86), .B1(new_n571), .B2(new_n207), .ZN(new_n573));
  NOR3_X1   g0373(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n257), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n385), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n545), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n385), .A2(new_n255), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n311), .A2(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n280), .A3(new_n282), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT85), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G116), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n280), .A3(new_n282), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n286), .ZN(new_n589));
  INV_X1    g0389(.A(G250), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n507), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n206), .A2(new_n293), .A3(G45), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n310), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G169), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n593), .ZN(new_n595));
  AOI211_X1 g0395(.A(G179), .B(new_n595), .C1(new_n588), .C2(new_n286), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n589), .A2(new_n451), .A3(new_n593), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n588), .B2(new_n286), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(G200), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n545), .A2(G87), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n576), .A2(new_n601), .A3(new_n579), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n580), .A2(new_n597), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n566), .A2(new_n567), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT89), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(G33), .B2(G283), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(G33), .B2(new_n284), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  AOI22_X1  g0410(.A1(KEYINPUT88), .A2(new_n609), .B1(new_n610), .B2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n611), .A3(new_n257), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n609), .A2(KEYINPUT88), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n255), .A2(G116), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n258), .B1(G1), .B2(new_n262), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(G116), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n308), .A2(G257), .A3(new_n345), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n308), .A2(G264), .A3(G1698), .ZN(new_n620));
  INV_X1    g0420(.A(G303), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n308), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n286), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n514), .A2(G270), .A3(new_n310), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n518), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT87), .B1(new_n624), .B2(new_n518), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n618), .B1(new_n627), .B2(new_n451), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n518), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n518), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n370), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n606), .B1(new_n628), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(G190), .A3(new_n623), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT89), .A4(new_n618), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT25), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n252), .B2(G107), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n549), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n545), .A2(G107), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n280), .A2(new_n282), .A3(new_n207), .A4(G87), .ZN(new_n645));
  AND2_X1   g0445(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n646));
  NOR2_X1   g0446(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n308), .A2(new_n207), .A3(G87), .A4(new_n646), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n584), .A2(G20), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT23), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n207), .B2(G107), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n549), .A2(KEYINPUT23), .A3(G20), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n649), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT24), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT24), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n649), .A2(new_n650), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n644), .B1(new_n660), .B2(new_n257), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n590), .A2(G1698), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n280), .A3(new_n282), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(KEYINPUT92), .B(G294), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G33), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(G1698), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n662), .A2(new_n280), .A3(new_n282), .A4(KEYINPUT91), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n665), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n286), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT93), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n517), .A2(new_n296), .A3(new_n511), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(G264), .B2(new_n529), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(KEYINPUT93), .A3(new_n286), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G169), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n286), .A2(new_n670), .B1(new_n529), .B2(G264), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(G179), .A3(new_n518), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n661), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n660), .A2(new_n257), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n643), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n673), .A2(new_n675), .A3(new_n451), .A4(new_n676), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n529), .A2(G264), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n370), .B1(new_n686), .B2(new_n674), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT21), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n631), .A2(new_n632), .B1(new_n286), .B2(new_n622), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n612), .B(new_n613), .Z(new_n692));
  INV_X1    g0492(.A(new_n615), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n545), .B2(new_n610), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G169), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n690), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n414), .B1(new_n622), .B2(new_n286), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n631), .B2(new_n632), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n627), .A2(KEYINPUT21), .A3(G169), .A4(new_n695), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n639), .A2(new_n689), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n504), .A2(new_n605), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT94), .Z(G372));
  NOR2_X1   g0506(.A1(new_n417), .A2(new_n488), .ZN(new_n707));
  INV_X1    g0507(.A(new_n327), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n491), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT80), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n489), .A2(new_n249), .A3(new_n491), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n558), .A2(new_n562), .A3(new_n561), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n548), .A2(new_n555), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n603), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n599), .A2(G200), .ZN(new_n717));
  AOI211_X1 g0517(.A(G190), .B(new_n595), .C1(new_n588), .C2(new_n286), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n602), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n599), .A2(new_n414), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(new_n580), .C1(G169), .C2(new_n599), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT26), .B1(new_n722), .B2(new_n563), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(new_n723), .A3(new_n721), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n716), .A2(new_n723), .A3(new_n726), .A4(new_n721), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n684), .A2(new_n687), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n661), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n603), .A2(new_n729), .A3(new_n563), .A4(new_n556), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n678), .A2(new_n680), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n683), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n697), .A3(new_n701), .A4(new_n702), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n725), .A2(new_n727), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n712), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n493), .A2(new_n326), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(new_n323), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n461), .A2(new_n467), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT96), .B1(new_n442), .B2(new_n465), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT96), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n483), .A2(new_n742), .A3(new_n484), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT18), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT18), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n739), .A2(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n368), .B1(new_n747), .B2(new_n365), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n737), .A2(new_n748), .ZN(G369));
  NAND2_X1  g0549(.A1(new_n251), .A2(new_n207), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT27), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT27), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(new_n752), .A3(G213), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G343), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n733), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT97), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n661), .A2(new_n755), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n681), .A2(new_n688), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n681), .A2(new_n756), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n758), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n733), .A2(new_n729), .ZN(new_n764));
  OAI211_X1 g0564(.A(KEYINPUT97), .B(new_n761), .C1(new_n764), .C2(new_n759), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n703), .A2(new_n756), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G330), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n639), .B(new_n703), .C1(new_n618), .C2(new_n755), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n695), .A3(new_n756), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n766), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(G399));
  INV_X1    g0575(.A(new_n210), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G41), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n574), .A2(new_n610), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n777), .A2(new_n206), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(KEYINPUT98), .B1(new_n213), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(KEYINPUT98), .B2(new_n779), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  INV_X1    g0583(.A(KEYINPUT30), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n698), .B1(new_n625), .B2(new_n626), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n679), .A2(new_n531), .A3(new_n599), .A4(new_n532), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT99), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n589), .A2(new_n593), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(new_n789), .B1(new_n679), .B2(new_n518), .ZN(new_n790));
  AOI21_X1  g0590(.A(G179), .B1(new_n531), .B2(new_n532), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n790), .A2(new_n627), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n785), .A2(new_n786), .A3(new_n784), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n787), .B(new_n793), .C1(new_n794), .C2(KEYINPUT100), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n533), .A2(new_n789), .A3(new_n686), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(KEYINPUT30), .A3(new_n700), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT100), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n756), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT31), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n798), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n803), .A2(new_n804), .A3(new_n787), .A4(new_n793), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(KEYINPUT31), .A3(new_n756), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n566), .A2(new_n567), .A3(new_n603), .A4(new_n755), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n802), .B(new_n806), .C1(new_n704), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G330), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n722), .A2(new_n563), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(new_n714), .B1(new_n580), .B2(new_n597), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n603), .A2(new_n713), .A3(new_n715), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT26), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n771), .A2(new_n681), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n811), .B(new_n813), .C1(new_n814), .C2(new_n730), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n755), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT29), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT29), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n736), .A2(new_n818), .A3(new_n755), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n809), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n783), .B1(new_n820), .B2(G1), .ZN(G364));
  NOR2_X1   g0621(.A1(new_n250), .A2(G20), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n206), .B1(new_n822), .B2(G45), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n777), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n773), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n770), .A2(new_n769), .A3(new_n772), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n770), .A2(new_n772), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n776), .A2(new_n283), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G355), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G116), .B2(new_n210), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n776), .A2(new_n308), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n288), .B2(new_n214), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n244), .A2(new_n288), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n215), .B1(G20), .B2(new_n412), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n833), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n825), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n207), .A2(G190), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n414), .A2(G200), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n207), .A2(new_n414), .A3(new_n370), .A4(G190), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(KEYINPUT33), .B(G317), .Z(new_n854));
  OAI221_X1 g0654(.A(new_n283), .B1(new_n850), .B2(new_n851), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(G179), .A2(G200), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n207), .B1(new_n856), .B2(G190), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n666), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n370), .A2(G179), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n847), .A2(new_n856), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n862), .B1(new_n864), .B2(G329), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n207), .A2(new_n451), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n860), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n621), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n866), .A2(new_n869), .A3(new_n848), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n866), .B2(new_n848), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(G322), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G326), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n207), .A2(new_n414), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(G190), .A3(G200), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT104), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n877), .B(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n859), .B(new_n874), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n877), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n881), .A2(G50), .B1(new_n849), .B2(new_n387), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n872), .B2(new_n330), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT103), .Z(new_n884));
  INV_X1    g0684(.A(G159), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n863), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT32), .ZN(new_n887));
  INV_X1    g0687(.A(G87), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n308), .B1(new_n867), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G107), .B2(new_n862), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n857), .A2(new_n284), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(G68), .B2(new_n852), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n880), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n846), .B1(new_n894), .B2(new_n843), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n826), .A2(new_n828), .B1(new_n834), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G396));
  AOI22_X1  g0697(.A1(new_n724), .A2(KEYINPUT95), .B1(new_n731), .B2(new_n734), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n756), .B1(new_n898), .B2(new_n727), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n398), .A2(new_n756), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n493), .B1(new_n410), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n416), .A2(new_n756), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n899), .B(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n825), .B1(new_n904), .B2(new_n809), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n809), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n843), .A2(new_n829), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n825), .B1(new_n908), .B2(G77), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT106), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n283), .B1(new_n864), .B2(G132), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n330), .B2(new_n857), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n867), .A2(new_n219), .B1(new_n861), .B2(new_n259), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(KEYINPUT108), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(KEYINPUT108), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT34), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n881), .A2(G137), .B1(new_n849), .B2(G159), .ZN(new_n917));
  XNOR2_X1  g0717(.A(KEYINPUT107), .B(G143), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n917), .B1(new_n335), .B2(new_n853), .C1(new_n872), .C2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n916), .ZN(new_n921));
  INV_X1    g0721(.A(G283), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n853), .A2(new_n922), .B1(new_n877), .B2(new_n621), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n283), .B1(new_n867), .B2(new_n549), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n923), .A2(new_n891), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(G87), .A2(new_n862), .B1(new_n864), .B2(G311), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n610), .B2(new_n850), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G294), .B2(new_n873), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n920), .A2(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n843), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n910), .B1(new_n929), .B2(new_n930), .C1(new_n903), .C2(new_n830), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n906), .A2(new_n931), .ZN(G384));
  OR2_X1    g0732(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(G116), .A3(new_n216), .A4(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT36), .Z(new_n936));
  OAI211_X1 g0736(.A(new_n387), .B(new_n214), .C1(new_n330), .C2(new_n259), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n219), .A2(G68), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n206), .B(G13), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n741), .A2(new_n743), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT18), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n740), .B1(new_n944), .B2(new_n744), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n483), .A2(new_n754), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT37), .B1(new_n483), .B2(new_n484), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n459), .A3(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT37), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n459), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n952), .B2(new_n942), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n945), .A2(new_n946), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT38), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n259), .B1(new_n439), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT109), .B1(new_n958), .B2(new_n426), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT109), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n960), .B(new_n469), .C1(new_n472), .C2(new_n259), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n961), .A3(new_n432), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n421), .B1(new_n962), .B2(new_n431), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n459), .B1(new_n753), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n465), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT37), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n948), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n962), .A2(new_n431), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n468), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n754), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n488), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n967), .A2(KEYINPUT38), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n941), .B1(new_n956), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n323), .A2(new_n326), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n275), .A2(new_n756), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n323), .A2(new_n326), .A3(new_n976), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n902), .B(new_n901), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n808), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n969), .A2(new_n484), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n970), .A3(new_n459), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n983), .A2(KEYINPUT37), .B1(new_n952), .B2(new_n947), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n970), .B1(new_n500), .B2(new_n497), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n955), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n973), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(new_n808), .A3(new_n980), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n974), .A2(new_n981), .B1(new_n988), .B2(new_n941), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n712), .A2(new_n808), .ZN(new_n991));
  OAI21_X1  g0791(.A(G330), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n736), .A2(new_n755), .A3(new_n903), .ZN(new_n994));
  INV_X1    g0794(.A(new_n902), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n978), .A2(new_n979), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n987), .A3(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n323), .A2(new_n756), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n986), .A2(KEYINPUT39), .A3(new_n973), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n967), .A2(KEYINPUT38), .A3(new_n972), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n955), .B2(new_n954), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1001), .C1(new_n1003), .C2(KEYINPUT39), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n944), .A2(new_n744), .A3(new_n753), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n998), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n748), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n819), .A2(new_n817), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n712), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1006), .B(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n993), .A2(new_n1010), .B1(new_n206), .B2(new_n822), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n993), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n940), .B1(new_n1011), .B2(new_n1012), .ZN(G367));
  OAI21_X1  g0813(.A(new_n603), .B1(new_n602), .B2(new_n755), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n721), .A2(new_n602), .A3(new_n755), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1016), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT43), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n766), .A2(new_n767), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n757), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n715), .A2(new_n756), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1024), .A2(new_n563), .A3(new_n556), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n713), .A2(new_n715), .A3(new_n756), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(KEYINPUT42), .B2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n563), .A2(new_n756), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n766), .A2(new_n767), .A3(new_n1027), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT42), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1017), .B(new_n1020), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1033), .A3(new_n1019), .A4(new_n1018), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n774), .A2(new_n1028), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n777), .B(KEYINPUT41), .Z(new_n1042));
  INV_X1    g0842(.A(KEYINPUT45), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n1027), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1023), .A2(KEYINPUT44), .A3(new_n1028), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT44), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n768), .B2(new_n1027), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n774), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1046), .A2(new_n1050), .A3(new_n774), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n766), .A2(new_n767), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n1021), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n1055), .B2(new_n1021), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n818), .B1(new_n815), .B2(new_n755), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n899), .B2(new_n818), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n809), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1058), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1053), .A2(new_n1054), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1042), .B1(new_n1066), .B2(new_n820), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1041), .B1(new_n1067), .B2(new_n824), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n844), .B1(new_n210), .B2(new_n385), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n839), .A2(new_n240), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n825), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n283), .B1(new_n861), .B2(new_n284), .ZN(new_n1072));
  INV_X1    g0872(.A(G317), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n850), .A2(new_n922), .B1(new_n863), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(G107), .C2(new_n858), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n621), .B2(new_n872), .C1(new_n851), .C2(new_n879), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n867), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n852), .A2(new_n666), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT46), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n867), .B2(new_n610), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT111), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n867), .A2(new_n330), .B1(new_n861), .B2(new_n226), .ZN(new_n1084));
  INV_X1    g0884(.A(G137), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n308), .B1(new_n863), .B2(new_n1085), .C1(new_n853), .C2(new_n885), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G50), .C2(new_n849), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n879), .B2(new_n918), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n857), .A2(new_n259), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n873), .B2(G150), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT112), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n1076), .A2(new_n1083), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT47), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1071), .B1(new_n1093), .B2(new_n843), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1018), .A2(new_n833), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1068), .A2(new_n1096), .ZN(G387));
  NOR2_X1   g0897(.A1(new_n1065), .A2(new_n780), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n820), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n766), .A2(new_n832), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n835), .A2(new_n778), .B1(new_n549), .B2(new_n776), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n237), .A2(new_n288), .ZN(new_n1103));
  AOI211_X1 g0903(.A(G45), .B(new_n778), .C1(G68), .C2(G77), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT50), .B1(new_n388), .B2(new_n219), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n388), .A2(KEYINPUT50), .A3(new_n219), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n838), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1102), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n844), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n825), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n387), .A2(new_n1077), .B1(new_n864), .B2(G150), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n259), .B2(new_n850), .C1(new_n872), .C2(new_n219), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n308), .B1(new_n861), .B2(new_n284), .C1(new_n877), .C2(new_n885), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n853), .A2(new_n418), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n857), .A2(new_n385), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT113), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n308), .B1(new_n864), .B2(G326), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1077), .A2(new_n666), .B1(new_n858), .B2(G283), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G311), .A2(new_n852), .B1(new_n849), .B2(G303), .ZN(new_n1121));
  INV_X1    g0921(.A(G322), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n872), .B2(new_n1073), .C1(new_n879), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT48), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT114), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT115), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT49), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1119), .B1(new_n610), .B2(new_n861), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1118), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1101), .B(new_n1111), .C1(new_n1133), .C2(new_n843), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1099), .B2(new_n824), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1100), .A2(new_n1135), .ZN(G393));
  AND3_X1   g0936(.A1(new_n1046), .A2(new_n1050), .A3(new_n774), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n774), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1028), .A2(new_n833), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n844), .B1(new_n284), .B2(new_n210), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n839), .A2(new_n247), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n825), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n849), .A2(new_n388), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n259), .B2(new_n867), .C1(new_n863), .C2(new_n918), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n308), .B1(new_n861), .B2(new_n888), .C1(new_n853), .C2(new_n219), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n857), .A2(new_n202), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n873), .A2(G159), .B1(G150), .B2(new_n881), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT51), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT116), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n283), .B1(new_n861), .B2(new_n549), .C1(new_n853), .C2(new_n621), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G322), .A2(new_n864), .B1(new_n849), .B2(G294), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n922), .B2(new_n867), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G116), .C2(new_n858), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n872), .A2(new_n851), .B1(new_n1073), .B2(new_n877), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1155), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1143), .B1(new_n1166), .B2(new_n843), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1139), .A2(new_n824), .B1(new_n1140), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1060), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1056), .B1(new_n1057), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n820), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n1066), .A3(new_n777), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1168), .A2(new_n1173), .ZN(G390));
  OAI211_X1 g0974(.A(G330), .B(new_n808), .C1(new_n492), .C2(new_n503), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n748), .C1(new_n1063), .C2(new_n504), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT118), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT118), .B1(new_n1009), .B2(new_n1175), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1001), .B1(new_n1003), .B2(KEYINPUT39), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n997), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n994), .B2(new_n995), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1183), .B2(new_n1000), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n500), .B1(new_n745), .B2(new_n746), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n946), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n942), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT37), .B1(new_n1187), .B2(new_n951), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1185), .A2(new_n1186), .B1(new_n1188), .B2(new_n948), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n973), .B1(new_n1189), .B2(KEYINPUT38), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n816), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n901), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n902), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n999), .B(new_n1190), .C1(new_n1193), .C2(new_n1182), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1184), .A2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n808), .A2(G330), .A3(new_n903), .A4(new_n997), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1184), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n802), .A2(new_n806), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n807), .A2(new_n704), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G330), .B(new_n903), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1182), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1196), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1180), .A2(new_n1198), .A3(new_n1199), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1009), .A2(KEYINPUT118), .A3(new_n1175), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1203), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1206), .B1(new_n1203), .B2(new_n1196), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1184), .A2(new_n1196), .A3(new_n1194), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1196), .B1(new_n1184), .B2(new_n1194), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1211), .A2(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1208), .A2(new_n1217), .A3(new_n777), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1198), .A2(new_n824), .A3(new_n1199), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1181), .A2(new_n829), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n825), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n308), .B1(new_n861), .B2(new_n219), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT54), .B(G143), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n850), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G125), .C2(new_n864), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n867), .A2(new_n335), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT53), .ZN(new_n1227));
  INV_X1    g1027(.A(G128), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1226), .A2(new_n1227), .B1(new_n1228), .B2(new_n877), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1227), .B2(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n873), .A2(G132), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G137), .A2(new_n852), .B1(new_n858), .B2(G159), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n850), .A2(new_n284), .B1(new_n259), .B2(new_n861), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G294), .B2(new_n864), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n308), .B(new_n1147), .C1(G87), .C2(new_n1077), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n873), .A2(G116), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n881), .A2(G283), .B1(new_n852), .B2(G107), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n930), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n908), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1221), .B(new_n1240), .C1(new_n418), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1219), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1218), .A2(new_n1245), .ZN(G378));
  NAND2_X1  g1046(.A1(new_n754), .A2(new_n338), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n501), .B(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1248), .B(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n989), .B2(G330), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n988), .A2(new_n941), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1190), .A2(KEYINPUT40), .A3(new_n808), .A4(new_n980), .ZN(new_n1254));
  AND4_X1   g1054(.A1(G330), .A2(new_n1253), .A3(new_n1254), .A4(new_n1251), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1006), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(G330), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1250), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n998), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n989), .A2(G330), .A3(new_n1251), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(KEYINPUT120), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT120), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .A4(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n824), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1250), .A2(new_n829), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n825), .B1(new_n908), .B2(G50), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT119), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n308), .A2(G41), .ZN(new_n1269));
  AOI211_X1 g1069(.A(G50), .B(new_n1269), .C1(new_n262), .C2(new_n287), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G58), .A2(new_n862), .B1(new_n864), .B2(G283), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n385), .B2(new_n850), .C1(new_n872), .C2(new_n549), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n226), .B2(new_n867), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n853), .A2(new_n284), .B1(new_n877), .B2(new_n610), .ZN(new_n1274));
  OR4_X1    g1074(.A1(new_n1089), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT58), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1270), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n850), .A2(new_n1085), .B1(new_n867), .B2(new_n1223), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G132), .B2(new_n852), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n881), .A2(G125), .B1(new_n858), .B2(G150), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1279), .B(new_n1280), .C1(new_n1228), .C2(new_n872), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(KEYINPUT59), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(KEYINPUT59), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n262), .B(new_n287), .C1(new_n861), .C2(new_n885), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G124), .B2(new_n864), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1277), .B1(new_n1276), .B2(new_n1275), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1268), .B1(new_n1287), .B2(new_n843), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1266), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1265), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT57), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1211), .B1(new_n1293), .B2(new_n1207), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1291), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1208), .A2(new_n1180), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1291), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n780), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1290), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(G375));
  AND3_X1   g1100(.A1(new_n1211), .A2(KEYINPUT121), .A3(new_n1214), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT121), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1042), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1207), .A2(new_n824), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n825), .B1(new_n908), .B2(G68), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n308), .B(new_n1116), .C1(G107), .C2(new_n849), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n873), .A2(G283), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n881), .A2(G294), .B1(new_n852), .B2(G116), .ZN(new_n1311));
  OAI22_X1  g1111(.A1(new_n867), .A2(new_n284), .B1(new_n861), .B2(new_n202), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(G303), .B2(new_n864), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n873), .A2(G137), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n283), .B1(new_n862), .B2(G58), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(G159), .A2(new_n1077), .B1(new_n864), .B2(G128), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1223), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n881), .A2(G132), .B1(new_n852), .B2(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(G50), .A2(new_n858), .B1(new_n849), .B2(G150), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(KEYINPUT122), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1308), .B1(new_n1323), .B2(new_n843), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1324), .B1(new_n997), .B2(new_n830), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1307), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1306), .A2(new_n1327), .ZN(G381));
  NAND3_X1  g1128(.A1(new_n1100), .A2(new_n1135), .A3(new_n896), .ZN(new_n1329));
  NOR4_X1   g1129(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n780), .B1(new_n1331), .B2(new_n1305), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1244), .B1(new_n1332), .B2(new_n1208), .ZN(new_n1333));
  INV_X1    g1133(.A(G381), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1330), .A2(new_n1333), .A3(new_n1299), .A4(new_n1334), .ZN(G407));
  INV_X1    g1135(.A(G213), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(G343), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1299), .A2(new_n1333), .A3(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(G407), .A2(G213), .A3(new_n1338), .ZN(G409));
  NAND2_X1  g1139(.A1(G393), .A2(G396), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1329), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1068), .A2(new_n1096), .A3(G390), .ZN(new_n1342));
  AOI21_X1  g1142(.A(G390), .B1(new_n1068), .B2(new_n1096), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1341), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(G390), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1137), .A2(new_n1138), .A3(new_n1171), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1304), .B1(new_n1347), .B2(new_n1064), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1348), .B2(new_n823), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1096), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1345), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1341), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1068), .A2(new_n1096), .A3(G390), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1344), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1337), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1214), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT121), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1211), .A2(KEYINPUT121), .A3(new_n1214), .ZN(new_n1360));
  OAI21_X1  g1160(.A(KEYINPUT60), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n780), .B1(new_n1363), .B2(KEYINPUT60), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1362), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(G384), .B1(new_n1365), .B2(new_n1327), .ZN(new_n1366));
  INV_X1    g1166(.A(G384), .ZN(new_n1367));
  AOI211_X1 g1167(.A(new_n1367), .B(new_n1326), .C1(new_n1362), .C2(new_n1364), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  AOI211_X1 g1169(.A(new_n1333), .B(new_n1290), .C1(new_n1295), .C2(new_n1298), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1296), .A2(new_n1304), .A3(new_n1264), .A4(new_n1262), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n823), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1372), .B1(new_n1266), .B2(new_n1288), .ZN(new_n1373));
  AOI21_X1  g1173(.A(G378), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1374));
  OAI211_X1 g1174(.A(new_n1356), .B(new_n1369), .C1(new_n1370), .C2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT123), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1374), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1378), .B1(G375), .B2(new_n1333), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1379), .A2(KEYINPUT123), .A3(new_n1356), .A4(new_n1369), .ZN(new_n1380));
  AOI21_X1  g1180(.A(KEYINPUT62), .B1(new_n1377), .B2(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1375), .A2(KEYINPUT62), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1337), .A2(G2897), .ZN(new_n1383));
  XOR2_X1   g1183(.A(new_n1383), .B(KEYINPUT125), .Z(new_n1384));
  NAND2_X1  g1184(.A1(new_n1337), .A2(KEYINPUT124), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1384), .B1(new_n1369), .B2(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT60), .ZN(new_n1387));
  OAI21_X1  g1187(.A(new_n777), .B1(new_n1357), .B2(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1388), .B1(new_n1303), .B2(new_n1361), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1367), .B1(new_n1389), .B2(new_n1326), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1365), .A2(G384), .A3(new_n1327), .ZN(new_n1391));
  AND4_X1   g1191(.A1(new_n1390), .A2(new_n1391), .A3(new_n1385), .A4(new_n1384), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1374), .B1(G378), .B2(new_n1299), .ZN(new_n1393));
  OAI22_X1  g1193(.A1(new_n1386), .A2(new_n1392), .B1(new_n1337), .B2(new_n1393), .ZN(new_n1394));
  INV_X1    g1194(.A(KEYINPUT61), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1382), .A2(new_n1394), .A3(new_n1395), .ZN(new_n1396));
  OAI21_X1  g1196(.A(new_n1355), .B1(new_n1381), .B2(new_n1396), .ZN(new_n1397));
  INV_X1    g1197(.A(KEYINPUT63), .ZN(new_n1398));
  NAND3_X1  g1198(.A1(new_n1377), .A2(new_n1380), .A3(new_n1398), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT126), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1400), .B1(new_n1386), .B2(new_n1392), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1379), .A2(new_n1356), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1390), .A2(new_n1391), .A3(new_n1385), .ZN(new_n1403));
  INV_X1    g1203(.A(new_n1384), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1403), .A2(new_n1404), .ZN(new_n1405));
  NAND3_X1  g1205(.A1(new_n1369), .A2(new_n1385), .A3(new_n1384), .ZN(new_n1406));
  NAND3_X1  g1206(.A1(new_n1405), .A2(new_n1406), .A3(KEYINPUT126), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1401), .A2(new_n1402), .A3(new_n1407), .ZN(new_n1408));
  OR2_X1    g1208(.A1(new_n1375), .A2(new_n1398), .ZN(new_n1409));
  NOR2_X1   g1209(.A1(new_n1355), .A2(KEYINPUT61), .ZN(new_n1410));
  NAND4_X1  g1210(.A1(new_n1399), .A2(new_n1408), .A3(new_n1409), .A4(new_n1410), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1397), .A2(new_n1411), .ZN(G405));
  AND3_X1   g1212(.A1(new_n1344), .A2(new_n1369), .A3(new_n1354), .ZN(new_n1413));
  AOI21_X1  g1213(.A(new_n1369), .B1(new_n1344), .B2(new_n1354), .ZN(new_n1414));
  OAI21_X1  g1214(.A(KEYINPUT127), .B1(new_n1413), .B2(new_n1414), .ZN(new_n1415));
  NAND2_X1  g1215(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1416));
  NAND2_X1  g1216(.A1(new_n1355), .A2(new_n1416), .ZN(new_n1417));
  INV_X1    g1217(.A(KEYINPUT127), .ZN(new_n1418));
  NAND3_X1  g1218(.A1(new_n1344), .A2(new_n1369), .A3(new_n1354), .ZN(new_n1419));
  NAND3_X1  g1219(.A1(new_n1417), .A2(new_n1418), .A3(new_n1419), .ZN(new_n1420));
  NOR2_X1   g1220(.A1(new_n1299), .A2(G378), .ZN(new_n1421));
  NOR2_X1   g1221(.A1(new_n1421), .A2(new_n1370), .ZN(new_n1422));
  AND3_X1   g1222(.A1(new_n1415), .A2(new_n1420), .A3(new_n1422), .ZN(new_n1423));
  AOI21_X1  g1223(.A(new_n1422), .B1(new_n1415), .B2(new_n1420), .ZN(new_n1424));
  NOR2_X1   g1224(.A1(new_n1423), .A2(new_n1424), .ZN(G402));
endmodule


