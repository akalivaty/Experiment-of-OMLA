

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734;

  NAND2_X2 U370 ( .A1(n642), .A2(n643), .ZN(n648) );
  XNOR2_X1 U371 ( .A(n391), .B(n390), .ZN(n471) );
  XNOR2_X1 U372 ( .A(n389), .B(KEYINPUT3), .ZN(n391) );
  INV_X1 U373 ( .A(n542), .ZN(n548) );
  XNOR2_X2 U374 ( .A(n351), .B(n352), .ZN(n668) );
  AND2_X1 U375 ( .A1(n373), .A2(n376), .ZN(n356) );
  NOR2_X1 U376 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U377 ( .A1(n503), .A2(n502), .ZN(n505) );
  XNOR2_X1 U378 ( .A(n546), .B(n545), .ZN(n733) );
  NOR2_X1 U379 ( .A1(n663), .A2(n664), .ZN(n531) );
  OR2_X1 U380 ( .A1(n607), .A2(G902), .ZN(n474) );
  AND2_X2 U381 ( .A1(n374), .A2(n598), .ZN(n695) );
  AND2_X2 U382 ( .A1(n374), .A2(n598), .ZN(n350) );
  NAND2_X1 U383 ( .A1(n356), .A2(n371), .ZN(n374) );
  NAND2_X1 U384 ( .A1(n496), .A2(n495), .ZN(n351) );
  XNOR2_X1 U385 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n352) );
  AND2_X1 U386 ( .A1(n491), .A2(n572), .ZN(n353) );
  BUF_X1 U387 ( .A(n416), .Z(n354) );
  XNOR2_X1 U388 ( .A(n387), .B(G122), .ZN(n416) );
  XOR2_X2 U389 ( .A(G125), .B(G146), .Z(n426) );
  XNOR2_X2 U390 ( .A(n454), .B(n453), .ZN(n720) );
  XNOR2_X1 U391 ( .A(n575), .B(n406), .ZN(n558) );
  NAND2_X1 U392 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n378) );
  NOR2_X1 U393 ( .A1(n594), .A2(n380), .ZN(n375) );
  XNOR2_X1 U394 ( .A(G137), .B(G131), .ZN(n452) );
  XNOR2_X1 U395 ( .A(n541), .B(KEYINPUT28), .ZN(n544) );
  INV_X1 U396 ( .A(n642), .ZN(n570) );
  XNOR2_X1 U397 ( .A(n425), .B(n424), .ZN(n517) );
  INV_X1 U398 ( .A(G478), .ZN(n423) );
  INV_X1 U399 ( .A(G953), .ZN(n706) );
  XNOR2_X1 U400 ( .A(n688), .B(KEYINPUT82), .ZN(n367) );
  XNOR2_X1 U401 ( .A(n369), .B(n368), .ZN(n687) );
  XNOR2_X1 U402 ( .A(n582), .B(n581), .ZN(n596) );
  AND2_X1 U403 ( .A1(n580), .A2(n355), .ZN(n582) );
  XNOR2_X1 U404 ( .A(G143), .B(G131), .ZN(n431) );
  XOR2_X1 U405 ( .A(G113), .B(G104), .Z(n434) );
  XNOR2_X1 U406 ( .A(G128), .B(G110), .ZN(n476) );
  XOR2_X1 U407 ( .A(G119), .B(G137), .Z(n478) );
  INV_X1 U408 ( .A(KEYINPUT64), .ZN(n397) );
  AND2_X1 U409 ( .A1(n382), .A2(n380), .ZN(n379) );
  NAND2_X1 U410 ( .A1(n363), .A2(n377), .ZN(n376) );
  NAND2_X1 U411 ( .A1(n381), .A2(n378), .ZN(n377) );
  XNOR2_X1 U412 ( .A(G107), .B(G101), .ZN(n458) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT78), .ZN(n393) );
  XOR2_X1 U414 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n394) );
  INV_X1 U415 ( .A(KEYINPUT81), .ZN(n368) );
  XNOR2_X1 U416 ( .A(n553), .B(n361), .ZN(n583) );
  XNOR2_X1 U417 ( .A(n364), .B(KEYINPUT84), .ZN(n575) );
  XNOR2_X1 U418 ( .A(n485), .B(KEYINPUT25), .ZN(n486) );
  AND2_X1 U419 ( .A1(n490), .A2(n572), .ZN(n523) );
  XOR2_X1 U420 ( .A(KEYINPUT5), .B(G116), .Z(n469) );
  XNOR2_X1 U421 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n545) );
  OR2_X1 U422 ( .A1(n676), .A2(n559), .ZN(n546) );
  INV_X1 U423 ( .A(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(G75) );
  INV_X1 U425 ( .A(KEYINPUT53), .ZN(n365) );
  NAND2_X1 U426 ( .A1(n367), .A2(n359), .ZN(n366) );
  NOR2_X1 U427 ( .A1(n639), .A2(n358), .ZN(n355) );
  INV_X1 U428 ( .A(KEYINPUT66), .ZN(n380) );
  AND2_X1 U429 ( .A1(n448), .A2(n643), .ZN(n357) );
  AND2_X1 U430 ( .A1(n579), .A2(KEYINPUT47), .ZN(n358) );
  AND2_X1 U431 ( .A1(n706), .A2(n680), .ZN(n359) );
  AND2_X1 U432 ( .A1(n405), .A2(G210), .ZN(n360) );
  XNOR2_X1 U433 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n361) );
  XNOR2_X1 U434 ( .A(KEYINPUT70), .B(KEYINPUT0), .ZN(n362) );
  INV_X1 U435 ( .A(n594), .ZN(n381) );
  OR2_X1 U436 ( .A1(n381), .A2(n380), .ZN(n363) );
  INV_X1 U437 ( .A(KEYINPUT2), .ZN(n382) );
  NAND2_X1 U438 ( .A1(n530), .A2(n659), .ZN(n364) );
  XNOR2_X2 U439 ( .A(n404), .B(n360), .ZN(n530) );
  NAND2_X1 U440 ( .A1(n705), .A2(n681), .ZN(n369) );
  XNOR2_X2 U441 ( .A(n529), .B(n528), .ZN(n705) );
  XNOR2_X2 U442 ( .A(G101), .B(G119), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n426), .B(n417), .ZN(n396) );
  XNOR2_X2 U444 ( .A(G143), .B(G128), .ZN(n417) );
  NOR2_X2 U445 ( .A1(n370), .A2(n668), .ZN(n497) );
  NOR2_X1 U446 ( .A1(n370), .A2(n654), .ZN(n513) );
  INV_X1 U447 ( .A(n506), .ZN(n370) );
  XNOR2_X2 U448 ( .A(n413), .B(n362), .ZN(n506) );
  NAND2_X1 U449 ( .A1(n372), .A2(n379), .ZN(n371) );
  INV_X1 U450 ( .A(n593), .ZN(n372) );
  NAND2_X1 U451 ( .A1(n593), .A2(n375), .ZN(n373) );
  XNOR2_X1 U452 ( .A(n354), .B(n415), .ZN(n422) );
  XNOR2_X2 U453 ( .A(KEYINPUT40), .B(n554), .ZN(n732) );
  AND2_X2 U454 ( .A1(n583), .A2(n634), .ZN(n554) );
  XNOR2_X2 U455 ( .A(G110), .B(G104), .ZN(n455) );
  XNOR2_X2 U456 ( .A(n397), .B(G953), .ZN(n722) );
  INV_X1 U457 ( .A(KEYINPUT44), .ZN(n504) );
  INV_X1 U458 ( .A(n685), .ZN(n598) );
  XNOR2_X1 U459 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U460 ( .A(n422), .B(n421), .ZN(n696) );
  XNOR2_X1 U461 ( .A(n423), .B(KEYINPUT101), .ZN(n424) );
  OR2_X1 U462 ( .A1(n722), .A2(G952), .ZN(n616) );
  XNOR2_X1 U463 ( .A(n455), .B(KEYINPUT16), .ZN(n388) );
  INV_X1 U464 ( .A(G107), .ZN(n383) );
  NAND2_X1 U465 ( .A1(G116), .A2(n383), .ZN(n386) );
  INV_X1 U466 ( .A(G116), .ZN(n384) );
  NAND2_X1 U467 ( .A1(n384), .A2(G107), .ZN(n385) );
  NAND2_X1 U468 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U469 ( .A(n388), .B(n416), .ZN(n392) );
  XNOR2_X1 U470 ( .A(G113), .B(KEYINPUT87), .ZN(n390) );
  XNOR2_X1 U471 ( .A(n392), .B(n471), .ZN(n714) );
  XNOR2_X1 U472 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U473 ( .A(n396), .B(n395), .ZN(n401) );
  XOR2_X1 U474 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n399) );
  NAND2_X1 U475 ( .A1(G224), .A2(n722), .ZN(n398) );
  XNOR2_X1 U476 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U477 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U478 ( .A(n714), .B(n402), .ZN(n612) );
  XNOR2_X1 U479 ( .A(G902), .B(KEYINPUT15), .ZN(n594) );
  NAND2_X1 U480 ( .A1(n612), .A2(n594), .ZN(n404) );
  INV_X1 U481 ( .A(G902), .ZN(n440) );
  INV_X1 U482 ( .A(G237), .ZN(n403) );
  NAND2_X1 U483 ( .A1(n440), .A2(n403), .ZN(n405) );
  NAND2_X1 U484 ( .A1(n405), .A2(G214), .ZN(n659) );
  XNOR2_X1 U485 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n406) );
  NAND2_X1 U486 ( .A1(G234), .A2(G237), .ZN(n407) );
  XNOR2_X1 U487 ( .A(n407), .B(KEYINPUT14), .ZN(n408) );
  XNOR2_X1 U488 ( .A(KEYINPUT76), .B(n408), .ZN(n410) );
  NAND2_X1 U489 ( .A1(n410), .A2(G902), .ZN(n409) );
  XNOR2_X1 U490 ( .A(n409), .B(KEYINPUT89), .ZN(n532) );
  NOR2_X1 U491 ( .A1(G898), .A2(n706), .ZN(n713) );
  AND2_X1 U492 ( .A1(n532), .A2(n713), .ZN(n411) );
  NAND2_X1 U493 ( .A1(G952), .A2(n410), .ZN(n675) );
  NOR2_X1 U494 ( .A1(n675), .A2(G953), .ZN(n535) );
  NOR2_X1 U495 ( .A1(n411), .A2(n535), .ZN(n412) );
  NOR2_X2 U496 ( .A1(n558), .A2(n412), .ZN(n413) );
  NAND2_X1 U497 ( .A1(n722), .A2(G234), .ZN(n414) );
  XOR2_X1 U498 ( .A(KEYINPUT8), .B(n414), .Z(n475) );
  NAND2_X1 U499 ( .A1(G217), .A2(n475), .ZN(n415) );
  XNOR2_X2 U500 ( .A(n417), .B(G134), .ZN(n454) );
  XOR2_X1 U501 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n419) );
  XNOR2_X1 U502 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n418) );
  XNOR2_X1 U503 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U504 ( .A(n454), .B(n420), .Z(n421) );
  NOR2_X1 U505 ( .A1(G902), .A2(n696), .ZN(n425) );
  XNOR2_X1 U506 ( .A(n426), .B(G140), .ZN(n427) );
  XNOR2_X1 U507 ( .A(n427), .B(KEYINPUT10), .ZN(n718) );
  XOR2_X1 U508 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n429) );
  XNOR2_X1 U509 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n428) );
  XNOR2_X1 U510 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U511 ( .A(n430), .B(KEYINPUT97), .Z(n432) );
  XNOR2_X1 U512 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U513 ( .A(n718), .B(n433), .Z(n439) );
  NOR2_X1 U514 ( .A1(G953), .A2(G237), .ZN(n467) );
  NAND2_X1 U515 ( .A1(G214), .A2(n467), .ZN(n435) );
  XNOR2_X1 U516 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U517 ( .A(KEYINPUT11), .B(G122), .Z(n436) );
  XNOR2_X1 U518 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U519 ( .A(n439), .B(n438), .ZN(n600) );
  NAND2_X1 U520 ( .A1(n600), .A2(n440), .ZN(n442) );
  XNOR2_X1 U521 ( .A(KEYINPUT13), .B(G475), .ZN(n441) );
  XNOR2_X1 U522 ( .A(n442), .B(n441), .ZN(n515) );
  NAND2_X1 U523 ( .A1(n517), .A2(n515), .ZN(n663) );
  INV_X1 U524 ( .A(n663), .ZN(n448) );
  XOR2_X1 U525 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n444) );
  NAND2_X1 U526 ( .A1(G234), .A2(n594), .ZN(n443) );
  XNOR2_X1 U527 ( .A(n444), .B(n443), .ZN(n484) );
  NAND2_X1 U528 ( .A1(n484), .A2(G221), .ZN(n447) );
  INV_X1 U529 ( .A(KEYINPUT92), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n445), .B(KEYINPUT21), .ZN(n446) );
  XNOR2_X1 U531 ( .A(n447), .B(n446), .ZN(n643) );
  NAND2_X1 U532 ( .A1(n506), .A2(n357), .ZN(n451) );
  INV_X1 U533 ( .A(KEYINPUT68), .ZN(n449) );
  XNOR2_X1 U534 ( .A(n449), .B(KEYINPUT22), .ZN(n450) );
  XNOR2_X1 U535 ( .A(n451), .B(n450), .ZN(n490) );
  XNOR2_X1 U536 ( .A(n452), .B(KEYINPUT4), .ZN(n453) );
  XNOR2_X1 U537 ( .A(n720), .B(G146), .ZN(n473) );
  INV_X1 U538 ( .A(n473), .ZN(n462) );
  NAND2_X1 U539 ( .A1(n722), .A2(G227), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U541 ( .A(KEYINPUT90), .B(G140), .ZN(n457) );
  XNOR2_X1 U542 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U543 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U544 ( .A(n462), .B(n461), .ZN(n691) );
  OR2_X2 U545 ( .A1(n691), .A2(G902), .ZN(n465) );
  INV_X1 U546 ( .A(KEYINPUT73), .ZN(n463) );
  XNOR2_X1 U547 ( .A(n463), .B(G469), .ZN(n464) );
  XNOR2_X2 U548 ( .A(n465), .B(n464), .ZN(n542) );
  XNOR2_X1 U549 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n466) );
  XNOR2_X2 U550 ( .A(n548), .B(n466), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n467), .A2(G210), .ZN(n468) );
  XNOR2_X1 U552 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U554 ( .A(n473), .B(n472), .ZN(n607) );
  XNOR2_X2 U555 ( .A(n474), .B(G472), .ZN(n646) );
  INV_X1 U556 ( .A(n646), .ZN(n539) );
  NAND2_X1 U557 ( .A1(n475), .A2(G221), .ZN(n481) );
  XOR2_X1 U558 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n477) );
  XNOR2_X1 U559 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U560 ( .A(n481), .B(n480), .ZN(n483) );
  INV_X1 U561 ( .A(n718), .ZN(n482) );
  XNOR2_X1 U562 ( .A(n483), .B(n482), .ZN(n701) );
  NOR2_X1 U563 ( .A1(n701), .A2(G902), .ZN(n487) );
  NAND2_X1 U564 ( .A1(G217), .A2(n484), .ZN(n485) );
  XNOR2_X2 U565 ( .A(n487), .B(n486), .ZN(n642) );
  NAND2_X1 U566 ( .A1(n539), .A2(n570), .ZN(n488) );
  NOR2_X1 U567 ( .A1(n495), .A2(n488), .ZN(n489) );
  NAND2_X1 U568 ( .A1(n490), .A2(n489), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(G110), .ZN(G12) );
  XNOR2_X1 U570 ( .A(n646), .B(KEYINPUT6), .ZN(n572) );
  INV_X1 U571 ( .A(n495), .ZN(n649) );
  NOR2_X1 U572 ( .A1(n649), .A2(n642), .ZN(n491) );
  NAND2_X1 U573 ( .A1(n353), .A2(n490), .ZN(n494) );
  XOR2_X1 U574 ( .A(KEYINPUT79), .B(KEYINPUT32), .Z(n492) );
  XNOR2_X1 U575 ( .A(n492), .B(KEYINPUT67), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n494), .B(n493), .ZN(n503) );
  XOR2_X1 U577 ( .A(G119), .B(n503), .Z(G21) );
  NOR2_X1 U578 ( .A1(n648), .A2(n572), .ZN(n496) );
  XNOR2_X1 U579 ( .A(n497), .B(KEYINPUT34), .ZN(n498) );
  NOR2_X1 U580 ( .A1(n517), .A2(n515), .ZN(n563) );
  NAND2_X1 U581 ( .A1(n498), .A2(n563), .ZN(n500) );
  XNOR2_X2 U582 ( .A(n500), .B(n499), .ZN(n620) );
  NAND2_X1 U583 ( .A1(n620), .A2(n501), .ZN(n502) );
  XNOR2_X1 U584 ( .A(n505), .B(n504), .ZN(n522) );
  BUF_X1 U585 ( .A(n506), .Z(n509) );
  INV_X1 U586 ( .A(n648), .ZN(n511) );
  NAND2_X1 U587 ( .A1(n542), .A2(n511), .ZN(n507) );
  NOR2_X1 U588 ( .A1(n507), .A2(n646), .ZN(n508) );
  NAND2_X1 U589 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U590 ( .A(KEYINPUT93), .B(n510), .ZN(n623) );
  NAND2_X1 U591 ( .A1(n646), .A2(n511), .ZN(n512) );
  OR2_X1 U592 ( .A1(n649), .A2(n512), .ZN(n654) );
  XOR2_X1 U593 ( .A(KEYINPUT31), .B(n513), .Z(n637) );
  NOR2_X1 U594 ( .A1(n623), .A2(n637), .ZN(n514) );
  XNOR2_X1 U595 ( .A(n514), .B(KEYINPUT94), .ZN(n520) );
  INV_X1 U596 ( .A(n515), .ZN(n516) );
  NOR2_X1 U597 ( .A1(n517), .A2(n516), .ZN(n636) );
  INV_X1 U598 ( .A(n636), .ZN(n519) );
  AND2_X1 U599 ( .A1(n517), .A2(n516), .ZN(n634) );
  INV_X1 U600 ( .A(n634), .ZN(n518) );
  NAND2_X1 U601 ( .A1(n519), .A2(n518), .ZN(n578) );
  INV_X1 U602 ( .A(n578), .ZN(n665) );
  NOR2_X1 U603 ( .A1(n520), .A2(n665), .ZN(n521) );
  NAND2_X1 U604 ( .A1(n523), .A2(n649), .ZN(n524) );
  XNOR2_X1 U605 ( .A(n524), .B(KEYINPUT83), .ZN(n525) );
  NAND2_X1 U606 ( .A1(n525), .A2(n642), .ZN(n526) );
  XNOR2_X1 U607 ( .A(n526), .B(KEYINPUT102), .ZN(n734) );
  NAND2_X1 U608 ( .A1(n527), .A2(n734), .ZN(n529) );
  XNOR2_X1 U609 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n528) );
  BUF_X1 U610 ( .A(n530), .Z(n562) );
  INV_X1 U611 ( .A(n562), .ZN(n589) );
  XNOR2_X1 U612 ( .A(n589), .B(KEYINPUT38), .ZN(n660) );
  NAND2_X1 U613 ( .A1(n660), .A2(n659), .ZN(n664) );
  XNOR2_X1 U614 ( .A(KEYINPUT41), .B(n531), .ZN(n676) );
  INV_X1 U615 ( .A(n722), .ZN(n533) );
  NAND2_X1 U616 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U617 ( .A1(G900), .A2(n534), .ZN(n536) );
  NOR2_X1 U618 ( .A1(n536), .A2(n535), .ZN(n547) );
  INV_X1 U619 ( .A(n643), .ZN(n537) );
  NOR2_X1 U620 ( .A1(n547), .A2(n537), .ZN(n569) );
  INV_X1 U621 ( .A(n569), .ZN(n538) );
  NOR2_X1 U622 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U623 ( .A1(n570), .A2(n540), .ZN(n541) );
  XNOR2_X1 U624 ( .A(n542), .B(KEYINPUT106), .ZN(n543) );
  NAND2_X1 U625 ( .A1(n544), .A2(n543), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U627 ( .A1(n646), .A2(n659), .ZN(n549) );
  XOR2_X1 U628 ( .A(KEYINPUT30), .B(n549), .Z(n550) );
  NAND2_X1 U629 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X2 U630 ( .A1(n552), .A2(n648), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n561), .A2(n660), .ZN(n553) );
  NOR2_X2 U632 ( .A1(n733), .A2(n732), .ZN(n555) );
  XNOR2_X1 U633 ( .A(n555), .B(KEYINPUT46), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT71), .B(KEYINPUT47), .ZN(n556) );
  NAND2_X1 U635 ( .A1(n556), .A2(n578), .ZN(n557) );
  XNOR2_X1 U636 ( .A(n557), .B(KEYINPUT75), .ZN(n560) );
  NOR2_X1 U637 ( .A1(n559), .A2(n558), .ZN(n632) );
  NAND2_X1 U638 ( .A1(n560), .A2(n632), .ZN(n566) );
  INV_X1 U639 ( .A(n561), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n563), .A2(n562), .ZN(n564) );
  OR2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n631) );
  AND2_X1 U642 ( .A1(n566), .A2(n631), .ZN(n567) );
  AND2_X1 U643 ( .A1(n568), .A2(n567), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U645 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U646 ( .A(n573), .B(KEYINPUT103), .Z(n574) );
  NAND2_X1 U647 ( .A1(n634), .A2(n574), .ZN(n584) );
  OR2_X1 U648 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U649 ( .A(n576), .B(KEYINPUT36), .ZN(n577) );
  NOR2_X1 U650 ( .A1(n577), .A2(n649), .ZN(n639) );
  NAND2_X1 U651 ( .A1(n632), .A2(n578), .ZN(n579) );
  XNOR2_X1 U652 ( .A(KEYINPUT48), .B(KEYINPUT72), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n636), .A2(n583), .ZN(n641) );
  INV_X1 U654 ( .A(n584), .ZN(n585) );
  AND2_X1 U655 ( .A1(n659), .A2(n585), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n649), .A2(n586), .ZN(n588) );
  XNOR2_X1 U657 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n588), .B(n587), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT105), .ZN(n730) );
  INV_X1 U661 ( .A(n730), .ZN(n592) );
  AND2_X1 U662 ( .A1(n641), .A2(n592), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n721) );
  NOR2_X2 U664 ( .A1(n705), .A2(n721), .ZN(n593) );
  AND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n683) );
  NAND2_X1 U666 ( .A1(n683), .A2(KEYINPUT2), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n705), .A2(n597), .ZN(n685) );
  NAND2_X1 U668 ( .A1(n350), .A2(G475), .ZN(n602) );
  XNOR2_X1 U669 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(n616), .ZN(n605) );
  XOR2_X1 U673 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(G60) );
  NAND2_X1 U675 ( .A1(n350), .A2(G472), .ZN(n609) );
  XOR2_X1 U676 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U678 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n610), .A2(n616), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n611), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U681 ( .A1(n695), .A2(G210), .ZN(n615) );
  XNOR2_X1 U682 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n612), .B(n613), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(n617) );
  INV_X1 U685 ( .A(n616), .ZN(n704) );
  NOR2_X2 U686 ( .A1(n617), .A2(n704), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n618), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U688 ( .A(G122), .B(KEYINPUT127), .Z(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(G24) );
  XOR2_X1 U690 ( .A(G104), .B(KEYINPUT109), .Z(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n634), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G6) );
  XNOR2_X1 U693 ( .A(G107), .B(KEYINPUT27), .ZN(n627) );
  XOR2_X1 U694 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n625) );
  NAND2_X1 U695 ( .A1(n623), .A2(n636), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(G9) );
  XOR2_X1 U698 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n629) );
  NAND2_X1 U699 ( .A1(n632), .A2(n636), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(G128), .B(n630), .Z(G30) );
  XNOR2_X1 U702 ( .A(G143), .B(n631), .ZN(G45) );
  NAND2_X1 U703 ( .A1(n632), .A2(n634), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(G146), .ZN(G48) );
  NAND2_X1 U705 ( .A1(n637), .A2(n634), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n635), .B(G113), .ZN(G15) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(G116), .ZN(G18) );
  XNOR2_X1 U709 ( .A(n639), .B(G125), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G134), .B(n641), .ZN(G36) );
  NOR2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U713 ( .A(KEYINPUT49), .B(n644), .Z(n645) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT113), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n650) );
  XNOR2_X1 U718 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n656) );
  INV_X1 U720 ( .A(n654), .ZN(n655) );
  NOR2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U722 ( .A(KEYINPUT51), .B(n657), .Z(n658) );
  NOR2_X1 U723 ( .A1(n676), .A2(n658), .ZN(n671) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT115), .B(n661), .Z(n662) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U730 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U731 ( .A(n672), .B(KEYINPUT52), .ZN(n673) );
  XNOR2_X1 U732 ( .A(KEYINPUT116), .B(n673), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n675), .A2(n674), .ZN(n678) );
  NOR2_X1 U734 ( .A1(n676), .A2(n668), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U736 ( .A(KEYINPUT117), .B(n679), .Z(n680) );
  XNOR2_X1 U737 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n682) );
  INV_X1 U738 ( .A(n682), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U740 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U741 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U742 ( .A1(n350), .A2(G469), .ZN(n693) );
  XNOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n689) );
  XOR2_X1 U744 ( .A(n689), .B(KEYINPUT57), .Z(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n704), .A2(n694), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n695), .A2(G478), .ZN(n698) );
  XOR2_X1 U749 ( .A(n696), .B(KEYINPUT121), .Z(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X2 U751 ( .A1(n699), .A2(n704), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n700), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U753 ( .A1(n350), .A2(G217), .ZN(n702) );
  XNOR2_X1 U754 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n704), .A2(n703), .ZN(G66) );
  INV_X1 U756 ( .A(n705), .ZN(n707) );
  NAND2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n712) );
  XOR2_X1 U758 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n709) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U761 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U762 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U765 ( .A(KEYINPUT124), .B(n717), .ZN(G69) );
  XNOR2_X1 U766 ( .A(n718), .B(KEYINPUT125), .ZN(n719) );
  XOR2_X1 U767 ( .A(n720), .B(n719), .Z(n725) );
  XNOR2_X1 U768 ( .A(n721), .B(n725), .ZN(n723) );
  NAND2_X1 U769 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U770 ( .A(n724), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U771 ( .A(n725), .B(G227), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U774 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U775 ( .A(G140), .B(n730), .Z(n731) );
  XNOR2_X1 U776 ( .A(KEYINPUT112), .B(n731), .ZN(G42) );
  XOR2_X1 U777 ( .A(G131), .B(n732), .Z(G33) );
  XOR2_X1 U778 ( .A(n733), .B(G137), .Z(G39) );
  XNOR2_X1 U779 ( .A(G101), .B(n734), .ZN(G3) );
endmodule

