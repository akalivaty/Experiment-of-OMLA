

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786;

  XNOR2_X1 U384 ( .A(n551), .B(n387), .ZN(n581) );
  XNOR2_X1 U385 ( .A(n447), .B(KEYINPUT8), .ZN(n508) );
  NAND2_X1 U386 ( .A1(n705), .A2(n672), .ZN(n663) );
  XNOR2_X2 U387 ( .A(n650), .B(KEYINPUT76), .ZN(n705) );
  XNOR2_X2 U388 ( .A(n393), .B(n507), .ZN(n560) );
  XNOR2_X2 U389 ( .A(n390), .B(n457), .ZN(n549) );
  INV_X2 U390 ( .A(KEYINPUT64), .ZN(n439) );
  XOR2_X1 U391 ( .A(n624), .B(KEYINPUT36), .Z(n363) );
  XNOR2_X2 U392 ( .A(n599), .B(n408), .ZN(n407) );
  XNOR2_X1 U393 ( .A(n404), .B(KEYINPUT45), .ZN(n649) );
  XNOR2_X1 U394 ( .A(n421), .B(KEYINPUT40), .ZN(n605) );
  XNOR2_X1 U395 ( .A(n394), .B(KEYINPUT77), .ZN(n506) );
  XNOR2_X1 U396 ( .A(n534), .B(n420), .ZN(n710) );
  XNOR2_X1 U397 ( .A(n518), .B(n517), .ZN(n563) );
  XNOR2_X1 U398 ( .A(n379), .B(n378), .ZN(n389) );
  XNOR2_X1 U399 ( .A(n381), .B(n380), .ZN(n379) );
  NOR2_X1 U400 ( .A1(n508), .A2(n509), .ZN(n512) );
  XNOR2_X1 U401 ( .A(G128), .B(G143), .ZN(n495) );
  BUF_X1 U402 ( .A(n428), .Z(n364) );
  NAND2_X1 U403 ( .A1(n364), .A2(n427), .ZN(n365) );
  NAND2_X1 U404 ( .A1(n428), .A2(n427), .ZN(n575) );
  BUF_X1 U405 ( .A(n571), .Z(n366) );
  XNOR2_X1 U406 ( .A(n415), .B(n369), .ZN(n535) );
  BUF_X1 U407 ( .A(n705), .Z(n367) );
  BUF_X1 U408 ( .A(n548), .Z(n368) );
  XNOR2_X2 U409 ( .A(n571), .B(KEYINPUT105), .ZN(n572) );
  NAND2_X2 U410 ( .A1(n565), .A2(n406), .ZN(n571) );
  XNOR2_X2 U411 ( .A(n576), .B(KEYINPUT87), .ZN(n403) );
  NOR2_X1 U412 ( .A1(n710), .A2(n418), .ZN(n712) );
  NAND2_X1 U413 ( .A1(n405), .A2(n407), .ZN(n397) );
  INV_X1 U414 ( .A(n719), .ZN(n405) );
  INV_X1 U415 ( .A(n718), .ZN(n547) );
  NAND2_X1 U416 ( .A1(n609), .A2(n372), .ZN(n433) );
  INV_X1 U417 ( .A(KEYINPUT78), .ZN(n423) );
  OR2_X1 U418 ( .A1(n666), .A2(G902), .ZN(n480) );
  NAND2_X1 U419 ( .A1(n448), .A2(G221), .ZN(n381) );
  XNOR2_X1 U420 ( .A(n454), .B(n451), .ZN(n380) );
  XNOR2_X1 U421 ( .A(G128), .B(G110), .ZN(n453) );
  XNOR2_X1 U422 ( .A(n510), .B(G122), .ZN(n511) );
  XNOR2_X1 U423 ( .A(n495), .B(n435), .ZN(n513) );
  XNOR2_X1 U424 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n449) );
  XNOR2_X1 U425 ( .A(n634), .B(n633), .ZN(n392) );
  XNOR2_X1 U426 ( .A(n417), .B(n377), .ZN(n739) );
  NOR2_X1 U427 ( .A1(n593), .A2(n594), .ZN(n417) );
  NAND2_X1 U428 ( .A1(n506), .A2(n419), .ZN(n393) );
  INV_X1 U429 ( .A(n710), .ZN(n419) );
  INV_X1 U430 ( .A(KEYINPUT1), .ZN(n408) );
  NAND2_X1 U431 ( .A1(n581), .A2(n386), .ZN(n554) );
  NAND2_X1 U432 ( .A1(n389), .A2(n388), .ZN(n390) );
  NOR2_X1 U433 ( .A1(n597), .A2(n573), .ZN(n431) );
  XNOR2_X1 U434 ( .A(n516), .B(KEYINPUT101), .ZN(n517) );
  BUF_X1 U435 ( .A(n492), .Z(n682) );
  XNOR2_X1 U436 ( .A(G902), .B(KEYINPUT15), .ZN(n642) );
  XOR2_X1 U437 ( .A(KEYINPUT5), .B(G146), .Z(n475) );
  XNOR2_X1 U438 ( .A(n513), .B(n436), .ZN(n474) );
  INV_X1 U439 ( .A(KEYINPUT44), .ZN(n411) );
  INV_X1 U440 ( .A(KEYINPUT38), .ZN(n420) );
  INV_X1 U441 ( .A(n619), .ZN(n386) );
  INV_X1 U442 ( .A(KEYINPUT74), .ZN(n387) );
  OR2_X1 U443 ( .A1(n700), .A2(G902), .ZN(n446) );
  XOR2_X1 U444 ( .A(G140), .B(G104), .Z(n524) );
  XNOR2_X1 U445 ( .A(n474), .B(n450), .ZN(n679) );
  INV_X1 U446 ( .A(G953), .ZN(n775) );
  AND2_X1 U447 ( .A1(n384), .A2(n375), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n385), .A2(n371), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n555), .A2(KEYINPUT34), .ZN(n410) );
  INV_X1 U450 ( .A(KEYINPUT22), .ZN(n412) );
  NOR2_X1 U451 ( .A1(n566), .A2(n396), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n397), .B(KEYINPUT104), .ZN(n396) );
  NAND2_X1 U453 ( .A1(n490), .A2(n489), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n424), .B(n423), .ZN(n490) );
  XNOR2_X1 U455 ( .A(n537), .B(n370), .ZN(n609) );
  XNOR2_X1 U456 ( .A(n549), .B(n398), .ZN(n719) );
  INV_X1 U457 ( .A(KEYINPUT103), .ZN(n398) );
  XNOR2_X1 U458 ( .A(G110), .B(G107), .ZN(n438) );
  XNOR2_X1 U459 ( .A(n678), .B(n452), .ZN(n378) );
  XNOR2_X1 U460 ( .A(n513), .B(n434), .ZN(n514) );
  XOR2_X1 U461 ( .A(G116), .B(G107), .Z(n434) );
  XNOR2_X1 U462 ( .A(n660), .B(KEYINPUT91), .ZN(n703) );
  NAND2_X1 U463 ( .A1(n392), .A2(n373), .ZN(n391) );
  INV_X1 U464 ( .A(G140), .ZN(n768) );
  XNOR2_X1 U465 ( .A(n416), .B(n603), .ZN(n786) );
  NAND2_X1 U466 ( .A1(n422), .A2(n564), .ZN(n421) );
  NAND2_X1 U467 ( .A1(n429), .A2(KEYINPUT66), .ZN(n427) );
  NOR2_X1 U468 ( .A1(n431), .A2(n549), .ZN(n430) );
  XOR2_X1 U469 ( .A(n505), .B(KEYINPUT92), .Z(n369) );
  XOR2_X1 U470 ( .A(n536), .B(KEYINPUT68), .Z(n370) );
  AND2_X1 U471 ( .A1(n368), .A2(n556), .ZN(n371) );
  XOR2_X1 U472 ( .A(n544), .B(KEYINPUT97), .Z(n372) );
  NAND2_X1 U473 ( .A1(n549), .A2(n718), .ZN(n721) );
  AND2_X1 U474 ( .A1(n639), .A2(KEYINPUT2), .ZN(n373) );
  AND2_X1 U475 ( .A1(n597), .A2(n573), .ZN(n374) );
  AND2_X1 U476 ( .A1(n410), .A2(n628), .ZN(n375) );
  XOR2_X1 U477 ( .A(n545), .B(KEYINPUT0), .Z(n376) );
  XNOR2_X1 U478 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n377) );
  XNOR2_X1 U479 ( .A(n485), .B(n484), .ZN(n709) );
  INV_X1 U480 ( .A(n709), .ZN(n418) );
  INV_X1 U481 ( .A(n389), .ZN(n690) );
  XNOR2_X2 U482 ( .A(n382), .B(n558), .ZN(n579) );
  NAND2_X1 U483 ( .A1(n383), .A2(n409), .ZN(n382) );
  INV_X1 U484 ( .A(n740), .ZN(n385) );
  INV_X1 U485 ( .A(G902), .ZN(n388) );
  AND2_X1 U486 ( .A1(n392), .A2(n639), .ZN(n647) );
  XNOR2_X1 U487 ( .A(n391), .B(KEYINPUT85), .ZN(n648) );
  XNOR2_X1 U488 ( .A(n395), .B(KEYINPUT80), .ZN(n567) );
  NAND2_X1 U489 ( .A1(n401), .A2(n399), .ZN(n404) );
  AND2_X1 U490 ( .A1(n400), .A2(n591), .ZN(n399) );
  NAND2_X1 U491 ( .A1(n580), .A2(n403), .ZN(n400) );
  XNOR2_X1 U492 ( .A(n402), .B(n411), .ZN(n401) );
  NAND2_X1 U493 ( .A1(n578), .A2(n403), .ZN(n402) );
  INV_X1 U494 ( .A(n407), .ZN(n406) );
  NAND2_X1 U495 ( .A1(n426), .A2(n407), .ZN(n551) );
  NAND2_X1 U496 ( .A1(n721), .A2(n406), .ZN(n722) );
  NAND2_X1 U497 ( .A1(n635), .A2(n406), .ZN(n636) );
  NAND2_X1 U498 ( .A1(n363), .A2(n407), .ZN(n767) );
  NAND2_X1 U499 ( .A1(n740), .A2(KEYINPUT34), .ZN(n409) );
  XNOR2_X2 U500 ( .A(n554), .B(n553), .ZN(n740) );
  XNOR2_X2 U501 ( .A(n413), .B(n412), .ZN(n565) );
  NAND2_X2 U502 ( .A1(n548), .A2(n414), .ZN(n413) );
  NOR2_X1 U503 ( .A1(n593), .A2(n547), .ZN(n414) );
  XNOR2_X2 U504 ( .A(n433), .B(n376), .ZN(n548) );
  INV_X1 U505 ( .A(n535), .ZN(n534) );
  NAND2_X1 U506 ( .A1(n652), .A2(n642), .ZN(n415) );
  XNOR2_X1 U507 ( .A(n503), .B(n771), .ZN(n652) );
  NAND2_X1 U508 ( .A1(n739), .A2(n608), .ZN(n416) );
  NAND2_X1 U509 ( .A1(n506), .A2(n623), .ZN(n627) );
  INV_X1 U510 ( .A(n605), .ZN(n592) );
  INV_X1 U511 ( .A(n560), .ZN(n422) );
  NAND2_X1 U512 ( .A1(n426), .A2(n425), .ZN(n424) );
  NOR2_X1 U513 ( .A1(n599), .A2(n595), .ZN(n425) );
  INV_X1 U514 ( .A(n721), .ZN(n426) );
  NAND2_X1 U515 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U516 ( .A(n572), .ZN(n429) );
  AND2_X2 U517 ( .A1(n432), .A2(n430), .ZN(n428) );
  NAND2_X1 U518 ( .A1(n572), .A2(n374), .ZN(n432) );
  INV_X1 U519 ( .A(n368), .ZN(n555) );
  AND2_X1 U520 ( .A1(n705), .A2(n672), .ZN(n689) );
  INV_X1 U521 ( .A(KEYINPUT66), .ZN(n573) );
  XNOR2_X1 U522 ( .A(n512), .B(n511), .ZN(n515) );
  INV_X1 U523 ( .A(G134), .ZN(n435) );
  XNOR2_X1 U524 ( .A(KEYINPUT4), .B(G131), .ZN(n436) );
  XNOR2_X1 U525 ( .A(n768), .B(G137), .ZN(n450) );
  INV_X1 U526 ( .A(G104), .ZN(n437) );
  XNOR2_X1 U527 ( .A(n438), .B(n437), .ZN(n772) );
  XNOR2_X1 U528 ( .A(n772), .B(KEYINPUT73), .ZN(n499) );
  XNOR2_X2 U529 ( .A(n439), .B(G953), .ZN(n492) );
  NAND2_X1 U530 ( .A1(n682), .A2(G227), .ZN(n441) );
  XOR2_X1 U531 ( .A(G146), .B(G101), .Z(n440) );
  XNOR2_X1 U532 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U533 ( .A(n499), .B(n442), .ZN(n443) );
  XNOR2_X1 U534 ( .A(n679), .B(n443), .ZN(n700) );
  INV_X1 U535 ( .A(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U536 ( .A(n444), .B(G469), .ZN(n445) );
  XNOR2_X2 U537 ( .A(n446), .B(n445), .ZN(n599) );
  NAND2_X1 U538 ( .A1(n492), .A2(G234), .ZN(n447) );
  INV_X1 U539 ( .A(n508), .ZN(n448) );
  INV_X1 U540 ( .A(G221), .ZN(n459) );
  XNOR2_X1 U541 ( .A(G146), .B(G125), .ZN(n496) );
  XNOR2_X1 U542 ( .A(n496), .B(n449), .ZN(n678) );
  INV_X1 U543 ( .A(n450), .ZN(n452) );
  XNOR2_X1 U544 ( .A(G119), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n453), .B(KEYINPUT23), .ZN(n454) );
  NAND2_X1 U546 ( .A1(n642), .A2(G234), .ZN(n455) );
  XNOR2_X1 U547 ( .A(n455), .B(KEYINPUT20), .ZN(n458) );
  AND2_X1 U548 ( .A1(n458), .A2(G217), .ZN(n456) );
  XNOR2_X1 U549 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  INV_X1 U550 ( .A(n458), .ZN(n460) );
  OR2_X1 U551 ( .A1(n460), .A2(n459), .ZN(n463) );
  INV_X1 U552 ( .A(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U553 ( .A(n461), .B(KEYINPUT21), .ZN(n462) );
  XNOR2_X1 U554 ( .A(n463), .B(n462), .ZN(n718) );
  NAND2_X1 U555 ( .A1(G234), .A2(G237), .ZN(n464) );
  XNOR2_X1 U556 ( .A(n464), .B(KEYINPUT94), .ZN(n465) );
  XNOR2_X1 U557 ( .A(KEYINPUT14), .B(n465), .ZN(n468) );
  AND2_X1 U558 ( .A1(n468), .A2(G952), .ZN(n736) );
  NAND2_X1 U559 ( .A1(n736), .A2(n775), .ZN(n467) );
  INV_X1 U560 ( .A(KEYINPUT95), .ZN(n466) );
  XNOR2_X1 U561 ( .A(n467), .B(n466), .ZN(n543) );
  NAND2_X1 U562 ( .A1(G902), .A2(n468), .ZN(n538) );
  NOR2_X1 U563 ( .A1(G900), .A2(n538), .ZN(n469) );
  INV_X1 U564 ( .A(n682), .ZN(n659) );
  NAND2_X1 U565 ( .A1(n469), .A2(n659), .ZN(n470) );
  AND2_X1 U566 ( .A1(n543), .A2(n470), .ZN(n595) );
  XNOR2_X1 U567 ( .A(G116), .B(G113), .ZN(n471) );
  XNOR2_X1 U568 ( .A(n471), .B(G119), .ZN(n473) );
  XNOR2_X1 U569 ( .A(G101), .B(KEYINPUT3), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n473), .B(n472), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n474), .B(n502), .ZN(n479) );
  NOR2_X1 U572 ( .A1(G953), .A2(G237), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n519), .A2(G210), .ZN(n477) );
  XNOR2_X1 U574 ( .A(n475), .B(G137), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n666) );
  XNOR2_X2 U577 ( .A(n480), .B(G472), .ZN(n727) );
  NOR2_X1 U578 ( .A1(G902), .A2(G237), .ZN(n482) );
  INV_X1 U579 ( .A(KEYINPUT75), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n482), .B(n481), .ZN(n504) );
  INV_X1 U581 ( .A(G214), .ZN(n483) );
  OR2_X1 U582 ( .A1(n504), .A2(n483), .ZN(n485) );
  INV_X1 U583 ( .A(KEYINPUT93), .ZN(n484) );
  NAND2_X1 U584 ( .A1(n727), .A2(n709), .ZN(n488) );
  XNOR2_X1 U585 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n486), .B(KEYINPUT108), .ZN(n487) );
  XNOR2_X1 U587 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X2 U588 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n491), .B(KEYINPUT4), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n492), .A2(G224), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n494), .B(n493), .ZN(n498) );
  XOR2_X1 U592 ( .A(n496), .B(n495), .Z(n497) );
  XNOR2_X1 U593 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U594 ( .A(n500), .B(n499), .ZN(n503) );
  XNOR2_X1 U595 ( .A(KEYINPUT16), .B(G122), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n771) );
  INV_X1 U597 ( .A(G210), .ZN(n651) );
  OR2_X1 U598 ( .A1(n504), .A2(n651), .ZN(n505) );
  INV_X1 U599 ( .A(KEYINPUT39), .ZN(n507) );
  INV_X1 U600 ( .A(G217), .ZN(n509) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n510) );
  XNOR2_X1 U602 ( .A(n515), .B(n514), .ZN(n693) );
  NOR2_X1 U603 ( .A1(G902), .A2(n693), .ZN(n518) );
  INV_X1 U604 ( .A(G478), .ZN(n516) );
  INV_X1 U605 ( .A(n563), .ZN(n533) );
  XOR2_X1 U606 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n521) );
  NAND2_X1 U607 ( .A1(G214), .A2(n519), .ZN(n520) );
  XNOR2_X1 U608 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U609 ( .A(n522), .B(n678), .Z(n530) );
  XNOR2_X1 U610 ( .A(G143), .B(G131), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n524), .B(n523), .ZN(n528) );
  XOR2_X1 U612 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n526) );
  XNOR2_X1 U613 ( .A(G113), .B(G122), .ZN(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U615 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n530), .B(n529), .ZN(n673) );
  NAND2_X1 U617 ( .A1(n673), .A2(n388), .ZN(n532) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(G475), .ZN(n531) );
  XNOR2_X1 U619 ( .A(n532), .B(n531), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n533), .A2(n561), .ZN(n764) );
  OR2_X1 U621 ( .A1(n560), .A2(n764), .ZN(n638) );
  XNOR2_X1 U622 ( .A(n638), .B(G134), .ZN(G36) );
  NAND2_X1 U623 ( .A1(n535), .A2(n709), .ZN(n537) );
  XNOR2_X1 U624 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n536) );
  INV_X1 U625 ( .A(n538), .ZN(n540) );
  INV_X1 U626 ( .A(G898), .ZN(n539) );
  AND2_X1 U627 ( .A1(n539), .A2(G953), .ZN(n773) );
  NAND2_X1 U628 ( .A1(n540), .A2(n773), .ZN(n541) );
  XNOR2_X1 U629 ( .A(n541), .B(KEYINPUT96), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n543), .A2(n542), .ZN(n544) );
  INV_X1 U631 ( .A(KEYINPUT69), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n563), .A2(n561), .ZN(n546) );
  XNOR2_X1 U633 ( .A(n546), .B(KEYINPUT102), .ZN(n593) );
  XNOR2_X1 U634 ( .A(n727), .B(KEYINPUT6), .ZN(n619) );
  NAND2_X1 U635 ( .A1(n619), .A2(n719), .ZN(n550) );
  NOR2_X1 U636 ( .A1(n366), .A2(n550), .ZN(n590) );
  XOR2_X1 U637 ( .A(G101), .B(n590), .Z(G3) );
  INV_X1 U638 ( .A(KEYINPUT90), .ZN(n552) );
  XNOR2_X1 U639 ( .A(n552), .B(KEYINPUT33), .ZN(n553) );
  INV_X1 U640 ( .A(KEYINPUT34), .ZN(n556) );
  NOR2_X1 U641 ( .A1(n563), .A2(n561), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT106), .ZN(n628) );
  XNOR2_X1 U643 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n558) );
  XNOR2_X1 U644 ( .A(G122), .B(KEYINPUT127), .ZN(n559) );
  XNOR2_X1 U645 ( .A(n579), .B(n559), .ZN(G24) );
  INV_X1 U646 ( .A(n561), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n761) );
  INV_X1 U648 ( .A(n761), .ZN(n564) );
  XOR2_X1 U649 ( .A(n592), .B(G131), .Z(G33) );
  XNOR2_X1 U650 ( .A(n619), .B(KEYINPUT81), .ZN(n566) );
  NAND2_X1 U651 ( .A1(n565), .A2(n567), .ZN(n570) );
  INV_X1 U652 ( .A(KEYINPUT65), .ZN(n568) );
  XNOR2_X1 U653 ( .A(n568), .B(KEYINPUT32), .ZN(n569) );
  XNOR2_X1 U654 ( .A(n570), .B(n569), .ZN(n574) );
  XNOR2_X1 U655 ( .A(n574), .B(G119), .ZN(G21) );
  INV_X1 U656 ( .A(n727), .ZN(n597) );
  XNOR2_X1 U657 ( .A(n365), .B(G110), .ZN(G12) );
  INV_X1 U658 ( .A(KEYINPUT70), .ZN(n577) );
  NOR2_X1 U659 ( .A1(n579), .A2(n577), .ZN(n578) );
  AND2_X1 U660 ( .A1(n579), .A2(n577), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n581), .A2(n727), .ZN(n729) );
  NOR2_X1 U662 ( .A1(n729), .A2(n555), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n582), .B(KEYINPUT31), .ZN(n763) );
  INV_X1 U664 ( .A(n763), .ZN(n586) );
  INV_X1 U665 ( .A(n599), .ZN(n584) );
  NOR2_X1 U666 ( .A1(n727), .A2(n721), .ZN(n583) );
  NAND2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U668 ( .A1(n555), .A2(n585), .ZN(n747) );
  NOR2_X1 U669 ( .A1(n586), .A2(n747), .ZN(n588) );
  AND2_X1 U670 ( .A1(n764), .A2(n761), .ZN(n612) );
  XOR2_X1 U671 ( .A(KEYINPUT83), .B(n612), .Z(n587) );
  NOR2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  BUF_X2 U674 ( .A(n649), .Z(n776) );
  INV_X1 U675 ( .A(n712), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n549), .A2(n595), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n596), .A2(n718), .ZN(n618) );
  NOR2_X1 U678 ( .A1(n618), .A2(n597), .ZN(n598) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(n598), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT111), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U682 ( .A(KEYINPUT112), .B(n602), .Z(n608) );
  INV_X1 U683 ( .A(KEYINPUT42), .ZN(n603) );
  INV_X1 U684 ( .A(n786), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U686 ( .A(KEYINPUT46), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n632) );
  AND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n759) );
  INV_X1 U689 ( .A(n612), .ZN(n711) );
  NAND2_X1 U690 ( .A1(n759), .A2(n711), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n610), .A2(KEYINPUT47), .ZN(n617) );
  NOR2_X1 U692 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n711), .A2(n611), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n612), .A2(KEYINPUT83), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n759), .A2(n615), .ZN(n616) );
  AND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n625) );
  OR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT107), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n621), .A2(n709), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n622), .A2(n761), .ZN(n635) );
  INV_X1 U702 ( .A(n534), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n635), .A2(n623), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n767), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT110), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n627), .B(n626), .ZN(n629) );
  AND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n757) );
  NOR2_X1 U708 ( .A1(n630), .A2(n757), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U710 ( .A(KEYINPUT48), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT43), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n637), .A2(n534), .ZN(n769) );
  AND2_X1 U713 ( .A1(n769), .A2(n638), .ZN(n639) );
  INV_X1 U714 ( .A(n647), .ZN(n640) );
  NOR2_X1 U715 ( .A1(n640), .A2(n642), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n776), .A2(n641), .ZN(n646) );
  XOR2_X1 U717 ( .A(KEYINPUT84), .B(n642), .Z(n643) );
  NAND2_X1 U718 ( .A1(n643), .A2(KEYINPUT2), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT67), .B(n644), .Z(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n672) );
  NAND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U722 ( .A1(n663), .A2(n651), .ZN(n657) );
  XNOR2_X1 U723 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n654) );
  XNOR2_X1 U724 ( .A(KEYINPUT55), .B(KEYINPUT82), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n652), .B(n655), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n661) );
  INV_X1 U728 ( .A(G952), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n703), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U732 ( .A(n663), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n664), .A2(G472), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U737 ( .A1(n669), .A2(n703), .ZN(n671) );
  XOR2_X1 U738 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G57) );
  NAND2_X1 U740 ( .A1(n689), .A2(G475), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT59), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X2 U743 ( .A1(n676), .A2(n703), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U745 ( .A(n679), .B(n678), .Z(n684) );
  INV_X1 U746 ( .A(n684), .ZN(n680) );
  XOR2_X1 U747 ( .A(KEYINPUT126), .B(n680), .Z(n681) );
  XNOR2_X1 U748 ( .A(n647), .B(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n688) );
  XOR2_X1 U750 ( .A(G227), .B(n684), .Z(n685) );
  NAND2_X1 U751 ( .A1(n685), .A2(G900), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n686), .A2(G953), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(G72) );
  BUF_X1 U754 ( .A(n689), .Z(n697) );
  NAND2_X1 U755 ( .A1(n697), .A2(G217), .ZN(n691) );
  XNOR2_X1 U756 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n692), .A2(n703), .ZN(G66) );
  NAND2_X1 U758 ( .A1(n697), .A2(G478), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT122), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n696), .A2(n703), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n697), .A2(G469), .ZN(n702) );
  XNOR2_X1 U763 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U764 ( .A(n698), .B(KEYINPUT58), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n776), .A2(n647), .ZN(n707) );
  INV_X1 U769 ( .A(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U771 ( .A1(n367), .A2(n708), .ZN(n745) );
  NAND2_X1 U772 ( .A1(n710), .A2(n418), .ZN(n715) );
  NAND2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U774 ( .A1(n593), .A2(n713), .ZN(n714) );
  NAND2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U776 ( .A1(n740), .A2(n716), .ZN(n717) );
  XOR2_X1 U777 ( .A(KEYINPUT120), .B(n717), .Z(n734) );
  NOR2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U779 ( .A(KEYINPUT49), .B(n720), .ZN(n725) );
  XNOR2_X1 U780 ( .A(n722), .B(KEYINPUT50), .ZN(n723) );
  XNOR2_X1 U781 ( .A(KEYINPUT118), .B(n723), .ZN(n724) );
  NAND2_X1 U782 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n728), .B(KEYINPUT119), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U786 ( .A(KEYINPUT51), .B(n731), .Z(n732) );
  NAND2_X1 U787 ( .A1(n739), .A2(n732), .ZN(n733) );
  NAND2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(KEYINPUT52), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n738), .A2(n775), .ZN(n743) );
  INV_X1 U792 ( .A(n739), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U796 ( .A(KEYINPUT53), .B(n746), .Z(G75) );
  INV_X1 U797 ( .A(n747), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n749), .A2(n761), .ZN(n748) );
  XOR2_X1 U799 ( .A(G104), .B(n748), .Z(G6) );
  NOR2_X1 U800 ( .A1(n749), .A2(n764), .ZN(n753) );
  XOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n751) );
  XNOR2_X1 U802 ( .A(G107), .B(KEYINPUT27), .ZN(n750) );
  XNOR2_X1 U803 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U804 ( .A(n753), .B(n752), .ZN(G9) );
  XOR2_X1 U805 ( .A(G128), .B(KEYINPUT29), .Z(n756) );
  INV_X1 U806 ( .A(n764), .ZN(n754) );
  NAND2_X1 U807 ( .A1(n759), .A2(n754), .ZN(n755) );
  XNOR2_X1 U808 ( .A(n756), .B(n755), .ZN(G30) );
  XOR2_X1 U809 ( .A(G143), .B(n757), .Z(n758) );
  XNOR2_X1 U810 ( .A(KEYINPUT116), .B(n758), .ZN(G45) );
  NAND2_X1 U811 ( .A1(n759), .A2(n564), .ZN(n760) );
  XNOR2_X1 U812 ( .A(G146), .B(n760), .ZN(G48) );
  NOR2_X1 U813 ( .A1(n761), .A2(n763), .ZN(n762) );
  XOR2_X1 U814 ( .A(G113), .B(n762), .Z(G15) );
  NOR2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U816 ( .A(G116), .B(n765), .Z(G18) );
  XOR2_X1 U817 ( .A(G125), .B(KEYINPUT37), .Z(n766) );
  XNOR2_X1 U818 ( .A(n767), .B(n766), .ZN(G27) );
  XNOR2_X1 U819 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U820 ( .A(n770), .B(KEYINPUT117), .ZN(G42) );
  XOR2_X1 U821 ( .A(n772), .B(n771), .Z(n774) );
  NOR2_X1 U822 ( .A1(n774), .A2(n773), .ZN(n785) );
  NAND2_X1 U823 ( .A1(n776), .A2(n775), .ZN(n782) );
  XOR2_X1 U824 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n778) );
  NAND2_X1 U825 ( .A1(G224), .A2(G953), .ZN(n777) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(n779) );
  NAND2_X1 U827 ( .A1(G898), .A2(n779), .ZN(n780) );
  XNOR2_X1 U828 ( .A(n780), .B(KEYINPUT124), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U830 ( .A(n783), .B(KEYINPUT125), .Z(n784) );
  XNOR2_X1 U831 ( .A(n785), .B(n784), .ZN(G69) );
  XOR2_X1 U832 ( .A(G137), .B(n786), .Z(G39) );
endmodule

