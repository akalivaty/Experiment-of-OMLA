

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588;

  INV_X1 U320 ( .A(KEYINPUT48), .ZN(n386) );
  XOR2_X1 U321 ( .A(n360), .B(KEYINPUT45), .Z(n288) );
  XOR2_X1 U322 ( .A(KEYINPUT70), .B(n324), .Z(n289) );
  NOR2_X1 U323 ( .A1(n382), .A2(n381), .ZN(n383) );
  INV_X1 U324 ( .A(G106GAT), .ZN(n333) );
  NOR2_X1 U325 ( .A1(n462), .A2(n538), .ZN(n388) );
  XNOR2_X1 U326 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U327 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U328 ( .A(n341), .B(n340), .ZN(n342) );
  NOR2_X1 U329 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U330 ( .A(n343), .B(n342), .ZN(n379) );
  XOR2_X1 U331 ( .A(n346), .B(n322), .Z(n579) );
  XNOR2_X1 U332 ( .A(n455), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n447), .B(G190GAT), .ZN(n448) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(G176GAT), .B(G204GAT), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n290), .B(G64GAT), .ZN(n319) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n323) );
  XOR2_X1 U338 ( .A(n319), .B(n323), .Z(n295) );
  XOR2_X1 U339 ( .A(G169GAT), .B(G8GAT), .Z(n363) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(KEYINPUT77), .Z(n292) );
  XNOR2_X1 U341 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U343 ( .A(KEYINPUT18), .B(n293), .Z(n444) );
  XNOR2_X1 U344 ( .A(n363), .B(n444), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U346 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n297) );
  NAND2_X1 U347 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(n299), .B(n298), .Z(n305) );
  XNOR2_X1 U350 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n300), .B(KEYINPUT80), .ZN(n301) );
  XOR2_X1 U352 ( .A(n301), .B(KEYINPUT81), .Z(n303) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n403) );
  XNOR2_X1 U355 ( .A(n403), .B(G92GAT), .ZN(n304) );
  XOR2_X1 U356 ( .A(n305), .B(n304), .Z(n526) );
  INV_X1 U357 ( .A(n526), .ZN(n462) );
  XNOR2_X1 U358 ( .A(G71GAT), .B(G57GAT), .ZN(n306) );
  XOR2_X1 U359 ( .A(n306), .B(KEYINPUT13), .Z(n346) );
  INV_X1 U360 ( .A(G92GAT), .ZN(n307) );
  NAND2_X1 U361 ( .A1(n307), .A2(KEYINPUT71), .ZN(n310) );
  INV_X1 U362 ( .A(KEYINPUT71), .ZN(n308) );
  NAND2_X1 U363 ( .A1(n308), .A2(G92GAT), .ZN(n309) );
  NAND2_X1 U364 ( .A1(n310), .A2(n309), .ZN(n312) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G85GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n324) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n289), .B(n313), .ZN(n317) );
  XOR2_X1 U369 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n315) );
  XNOR2_X1 U370 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U372 ( .A(n317), .B(n316), .Z(n321) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(G148GAT), .ZN(n402) );
  XNOR2_X1 U375 ( .A(n402), .B(n319), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  INV_X1 U377 ( .A(n579), .ZN(n475) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n328) );
  INV_X1 U379 ( .A(n328), .ZN(n326) );
  AND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  INV_X1 U381 ( .A(n327), .ZN(n325) );
  NAND2_X1 U382 ( .A1(n326), .A2(n325), .ZN(n330) );
  NAND2_X1 U383 ( .A1(n328), .A2(n327), .ZN(n329) );
  NAND2_X1 U384 ( .A1(n330), .A2(n329), .ZN(n336) );
  XOR2_X1 U385 ( .A(G29GAT), .B(G43GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n362) );
  XNOR2_X1 U388 ( .A(n362), .B(G134GAT), .ZN(n334) );
  XOR2_X1 U389 ( .A(n337), .B(KEYINPUT11), .Z(n343) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G162GAT), .Z(n391) );
  XNOR2_X1 U391 ( .A(G218GAT), .B(n391), .ZN(n341) );
  XOR2_X1 U392 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n339) );
  XNOR2_X1 U393 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(KEYINPUT36), .B(n379), .ZN(n491) );
  XOR2_X1 U396 ( .A(G155GAT), .B(G78GAT), .Z(n345) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n359) );
  XNOR2_X1 U399 ( .A(n346), .B(G127GAT), .ZN(n348) );
  XOR2_X1 U400 ( .A(G15GAT), .B(G1GAT), .Z(n374) );
  XNOR2_X1 U401 ( .A(n374), .B(G183GAT), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n350) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U406 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT12), .Z(n354) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(G64GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n355), .B(KEYINPUT74), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n458) );
  INV_X1 U413 ( .A(n458), .ZN(n572) );
  NOR2_X1 U414 ( .A1(n491), .A2(n572), .ZN(n360) );
  NOR2_X1 U415 ( .A1(n475), .A2(n288), .ZN(n361) );
  XNOR2_X1 U416 ( .A(KEYINPUT110), .B(n361), .ZN(n378) );
  XOR2_X1 U417 ( .A(G141GAT), .B(G22GAT), .Z(n392) );
  XNOR2_X1 U418 ( .A(n362), .B(n392), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n366) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n370) );
  XNOR2_X1 U425 ( .A(G113GAT), .B(G197GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT69), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U430 ( .A(G36GAT), .B(G50GAT), .ZN(n376) );
  XOR2_X1 U431 ( .A(n377), .B(n376), .Z(n505) );
  INV_X1 U432 ( .A(n505), .ZN(n574) );
  NAND2_X1 U433 ( .A1(n378), .A2(n574), .ZN(n385) );
  NAND2_X1 U434 ( .A1(n572), .A2(n379), .ZN(n382) );
  XOR2_X1 U435 ( .A(n579), .B(KEYINPUT41), .Z(n565) );
  NOR2_X1 U436 ( .A1(n574), .A2(n565), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n380), .B(KEYINPUT46), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n383), .B(KEYINPUT47), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n385), .A2(n384), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n538) );
  XNOR2_X1 U441 ( .A(n388), .B(KEYINPUT54), .ZN(n451) );
  XOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n390) );
  XNOR2_X1 U443 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n396) );
  XOR2_X1 U445 ( .A(G204GAT), .B(KEYINPUT84), .Z(n394) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U448 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n401) );
  XOR2_X1 U451 ( .A(G155GAT), .B(KEYINPUT82), .Z(n400) );
  XNOR2_X1 U452 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n420) );
  XOR2_X1 U454 ( .A(n401), .B(n420), .Z(n405) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n405), .B(n404), .ZN(n465) );
  XOR2_X1 U457 ( .A(G85GAT), .B(G148GAT), .Z(n407) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G141GAT), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U460 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n409) );
  XNOR2_X1 U461 ( .A(KEYINPUT1), .B(KEYINPUT86), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U463 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U464 ( .A(G127GAT), .B(G134GAT), .Z(n413) );
  XNOR2_X1 U465 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U467 ( .A(G113GAT), .B(n414), .Z(n438) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n416) );
  XNOR2_X1 U469 ( .A(G57GAT), .B(KEYINPUT85), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n438), .B(n417), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U473 ( .A(G162GAT), .B(n420), .Z(n422) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U476 ( .A(G29GAT), .B(n423), .Z(n424) );
  XOR2_X1 U477 ( .A(n425), .B(n424), .Z(n523) );
  NOR2_X1 U478 ( .A1(n465), .A2(n523), .ZN(n426) );
  AND2_X1 U479 ( .A1(n451), .A2(n426), .ZN(n428) );
  XNOR2_X1 U480 ( .A(KEYINPUT115), .B(KEYINPUT55), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n445) );
  XOR2_X1 U482 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n430) );
  XNOR2_X1 U483 ( .A(G15GAT), .B(G176GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT65), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G99GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U489 ( .A(G190GAT), .B(KEYINPUT76), .Z(n436) );
  XNOR2_X1 U490 ( .A(G43GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U492 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n463) );
  INV_X1 U497 ( .A(n463), .ZN(n540) );
  NAND2_X1 U498 ( .A1(n445), .A2(n540), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT116), .ZN(n571) );
  NOR2_X1 U500 ( .A1(n571), .A2(n379), .ZN(n449) );
  XNOR2_X1 U501 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n447) );
  INV_X1 U502 ( .A(G211GAT), .ZN(n457) );
  NAND2_X1 U503 ( .A1(n465), .A2(n463), .ZN(n450) );
  XOR2_X1 U504 ( .A(n450), .B(KEYINPUT26), .Z(n555) );
  INV_X1 U505 ( .A(n555), .ZN(n453) );
  INV_X1 U506 ( .A(n523), .ZN(n470) );
  NAND2_X1 U507 ( .A1(n451), .A2(n470), .ZN(n452) );
  XOR2_X1 U508 ( .A(KEYINPUT120), .B(n454), .Z(n586) );
  NOR2_X1 U509 ( .A1(n572), .A2(n586), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(G1354GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n479) );
  NAND2_X1 U512 ( .A1(n458), .A2(n379), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT75), .ZN(n474) );
  XNOR2_X1 U515 ( .A(n526), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U516 ( .A1(n523), .A2(n467), .ZN(n537) );
  NOR2_X1 U517 ( .A1(n540), .A2(n537), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n465), .B(KEYINPUT28), .ZN(n531) );
  INV_X1 U519 ( .A(n531), .ZN(n544) );
  NAND2_X1 U520 ( .A1(n461), .A2(n544), .ZN(n473) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n467), .A2(n555), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n489) );
  NAND2_X1 U528 ( .A1(n474), .A2(n489), .ZN(n507) );
  NOR2_X1 U529 ( .A1(n574), .A2(n475), .ZN(n476) );
  XOR2_X1 U530 ( .A(KEYINPUT72), .B(n476), .Z(n494) );
  NOR2_X1 U531 ( .A1(n507), .A2(n494), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT90), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n523), .A2(n486), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n486), .A2(n526), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT92), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT93), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U540 ( .A1(n486), .A2(n540), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(G15GAT), .B(n485), .Z(G1326GAT) );
  NAND2_X1 U543 ( .A1(n486), .A2(n531), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n487), .B(KEYINPUT94), .ZN(n488) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT95), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U547 ( .A1(n572), .A2(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT96), .B(n490), .ZN(n492) );
  NOR2_X1 U549 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(KEYINPUT37), .ZN(n521) );
  NOR2_X1 U551 ( .A1(n521), .A2(n494), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U553 ( .A1(n523), .A2(n503), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n498), .Z(G1328GAT) );
  NAND2_X1 U556 ( .A1(n503), .A2(n526), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT97), .Z(n501) );
  NAND2_X1 U559 ( .A1(n503), .A2(n540), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n531), .A2(n503), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT100), .B(KEYINPUT42), .Z(n510) );
  NOR2_X1 U565 ( .A1(n505), .A2(n565), .ZN(n506) );
  XOR2_X1 U566 ( .A(KEYINPUT98), .B(n506), .Z(n522) );
  NOR2_X1 U567 ( .A1(n522), .A2(n507), .ZN(n508) );
  XOR2_X1 U568 ( .A(KEYINPUT99), .B(n508), .Z(n516) );
  NAND2_X1 U569 ( .A1(n516), .A2(n523), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  XOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT101), .Z(n513) );
  NAND2_X1 U573 ( .A1(n516), .A2(n526), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n540), .A2(n516), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(KEYINPUT102), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U579 ( .A1(n516), .A2(n531), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT103), .Z(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT105), .Z(n525) );
  NOR2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n532), .A2(n523), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n532), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n527), .B(KEYINPUT106), .ZN(n528) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT107), .Z(n530) );
  NAND2_X1 U591 ( .A1(n532), .A2(n540), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n534) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(n536), .B(n535), .ZN(G1339GAT) );
  INV_X1 U598 ( .A(KEYINPUT112), .ZN(n542) );
  NOR2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT111), .B(n539), .Z(n556) );
  NAND2_X1 U601 ( .A1(n556), .A2(n540), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n551) );
  NOR2_X1 U604 ( .A1(n574), .A2(n551), .ZN(n545) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n545), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n565), .A2(n551), .ZN(n547) );
  XNOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  NOR2_X1 U610 ( .A1(n572), .A2(n551), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n379), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n562) );
  NOR2_X1 U618 ( .A1(n574), .A2(n562), .ZN(n557) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n557), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n565), .A2(n562), .ZN(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n572), .A2(n562), .ZN(n561) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n379), .A2(n562), .ZN(n563) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n574), .A2(n571), .ZN(n564) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n571), .A2(n565), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT118), .Z(n567) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT117), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT56), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  NOR2_X1 U638 ( .A1(n586), .A2(n574), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT121), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n586), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT123), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n491), .A2(n586), .ZN(n587) );
  XOR2_X1 U652 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

