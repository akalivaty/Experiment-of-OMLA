

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(n387), .B(n386), .ZN(n524) );
  NOR2_X1 U326 ( .A1(n389), .A2(n565), .ZN(n391) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n433) );
  XNOR2_X1 U328 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n466) );
  XNOR2_X1 U329 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U330 ( .A(G92GAT), .B(KEYINPUT68), .Z(n372) );
  INV_X1 U331 ( .A(KEYINPUT25), .ZN(n390) );
  XNOR2_X1 U332 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U333 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U334 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U335 ( .A(n444), .B(n443), .ZN(n465) );
  NOR2_X1 U336 ( .A1(n572), .A2(n571), .ZN(n580) );
  INV_X1 U337 ( .A(KEYINPUT112), .ZN(n462) );
  XOR2_X1 U338 ( .A(n420), .B(n419), .Z(n567) );
  XNOR2_X1 U339 ( .A(n462), .B(G50GAT), .ZN(n463) );
  XNOR2_X1 U340 ( .A(n464), .B(n463), .ZN(G1331GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n294) );
  XNOR2_X1 U342 ( .A(KEYINPUT94), .B(KEYINPUT89), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n311) );
  XOR2_X1 U344 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n296) );
  XNOR2_X1 U345 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U347 ( .A(n297), .B(KEYINPUT22), .Z(n299) );
  XOR2_X1 U348 ( .A(G141GAT), .B(G22GAT), .Z(n448) );
  XNOR2_X1 U349 ( .A(G50GAT), .B(n448), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U351 ( .A(G218GAT), .B(G162GAT), .Z(n322) );
  XOR2_X1 U352 ( .A(G211GAT), .B(KEYINPUT21), .Z(n301) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(KEYINPUT92), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n380) );
  XOR2_X1 U355 ( .A(n322), .B(n380), .Z(n303) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(n305), .B(n304), .Z(n309) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(G78GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U361 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n307), .B(KEYINPUT2), .ZN(n416) );
  XNOR2_X1 U363 ( .A(n439), .B(n416), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U365 ( .A(n311), .B(n310), .Z(n565) );
  XNOR2_X1 U366 ( .A(n565), .B(KEYINPUT28), .ZN(n537) );
  INV_X1 U367 ( .A(n537), .ZN(n528) );
  XOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT8), .Z(n313) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G36GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U371 ( .A(G50GAT), .B(KEYINPUT7), .Z(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n457) );
  INV_X1 U373 ( .A(n457), .ZN(n328) );
  XOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .Z(n434) );
  XOR2_X1 U375 ( .A(G134GAT), .B(KEYINPUT72), .Z(n400) );
  XOR2_X1 U376 ( .A(n434), .B(n400), .Z(n317) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U379 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n319) );
  XNOR2_X1 U380 ( .A(KEYINPUT73), .B(KEYINPUT9), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U382 ( .A(n321), .B(n320), .Z(n326) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n323), .B(G92GAT), .ZN(n324) );
  XNOR2_X1 U385 ( .A(G190GAT), .B(n324), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U387 ( .A(n328), .B(n327), .Z(n563) );
  XNOR2_X1 U388 ( .A(KEYINPUT36), .B(n563), .ZN(n483) );
  XOR2_X1 U389 ( .A(KEYINPUT74), .B(KEYINPUT77), .Z(n330) );
  XNOR2_X1 U390 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT13), .Z(n431) );
  XOR2_X1 U393 ( .A(n431), .B(G71GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G15GAT), .B(G1GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n331), .B(KEYINPUT66), .ZN(n447) );
  XNOR2_X1 U396 ( .A(n447), .B(G127GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n348) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G78GAT), .Z(n337) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U402 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n339) );
  XNOR2_X1 U403 ( .A(G211GAT), .B(G64GAT), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U405 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n343) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(n344), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n592) );
  INV_X1 U412 ( .A(n592), .ZN(n560) );
  XOR2_X1 U413 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT80), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U416 ( .A(G113GAT), .B(n351), .Z(n412) );
  XOR2_X1 U417 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n353) );
  XNOR2_X1 U418 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U420 ( .A(KEYINPUT88), .B(KEYINPUT82), .Z(n355) );
  XNOR2_X1 U421 ( .A(G169GAT), .B(G15GAT), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U423 ( .A(n357), .B(n356), .Z(n370) );
  XOR2_X1 U424 ( .A(G183GAT), .B(KEYINPUT85), .Z(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U427 ( .A(n360), .B(KEYINPUT17), .Z(n362) );
  XNOR2_X1 U428 ( .A(KEYINPUT19), .B(G190GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n387) );
  XOR2_X1 U430 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XOR2_X1 U431 ( .A(G176GAT), .B(G99GAT), .Z(n364) );
  XNOR2_X1 U432 ( .A(G43GAT), .B(G134GAT), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U434 ( .A(n440), .B(n365), .Z(n367) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n387), .B(n368), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n412), .B(n371), .ZN(n572) );
  XOR2_X1 U440 ( .A(G169GAT), .B(G8GAT), .Z(n451) );
  INV_X1 U441 ( .A(G204GAT), .ZN(n379) );
  XNOR2_X1 U442 ( .A(G176GAT), .B(G64GAT), .ZN(n373) );
  NAND2_X1 U443 ( .A1(n372), .A2(n373), .ZN(n377) );
  INV_X1 U444 ( .A(n372), .ZN(n375) );
  INV_X1 U445 ( .A(n373), .ZN(n374) );
  NAND2_X1 U446 ( .A1(n375), .A2(n374), .ZN(n376) );
  NAND2_X1 U447 ( .A1(n377), .A2(n376), .ZN(n378) );
  XOR2_X1 U448 ( .A(n433), .B(n380), .Z(n382) );
  XNOR2_X1 U449 ( .A(G36GAT), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U451 ( .A(n451), .B(n383), .Z(n385) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  NOR2_X1 U454 ( .A1(n572), .A2(n524), .ZN(n388) );
  XOR2_X1 U455 ( .A(KEYINPUT103), .B(n388), .Z(n389) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n395) );
  XNOR2_X1 U457 ( .A(KEYINPUT27), .B(n524), .ZN(n422) );
  NAND2_X1 U458 ( .A1(n572), .A2(n565), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT26), .ZN(n393) );
  XNOR2_X1 U460 ( .A(KEYINPUT102), .B(n393), .ZN(n480) );
  NOR2_X1 U461 ( .A1(n422), .A2(n480), .ZN(n394) );
  NOR2_X1 U462 ( .A1(n395), .A2(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(KEYINPUT104), .B(n396), .Z(n421) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G162GAT), .Z(n398) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G120GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U467 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n420) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n404) );
  XNOR2_X1 U471 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U473 ( .A(G57GAT), .B(G148GAT), .Z(n406) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(G1GAT), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U476 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U477 ( .A(KEYINPUT4), .B(KEYINPUT98), .Z(n410) );
  XNOR2_X1 U478 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U482 ( .A(n415), .B(KEYINPUT99), .Z(n418) );
  XNOR2_X1 U483 ( .A(n416), .B(KEYINPUT100), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U485 ( .A1(n421), .A2(n567), .ZN(n426) );
  NOR2_X1 U486 ( .A1(n422), .A2(n567), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n423), .B(KEYINPUT101), .ZN(n532) );
  NOR2_X1 U488 ( .A1(n537), .A2(n532), .ZN(n424) );
  NAND2_X1 U489 ( .A1(n424), .A2(n572), .ZN(n425) );
  NAND2_X1 U490 ( .A1(n426), .A2(n425), .ZN(n489) );
  NAND2_X1 U491 ( .A1(n560), .A2(n489), .ZN(n427) );
  NOR2_X1 U492 ( .A1(n483), .A2(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n521) );
  XOR2_X1 U495 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n430) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n444) );
  XOR2_X1 U497 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n437) );
  NAND2_X1 U498 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT31), .B(n438), .Z(n442) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(KEYINPUT30), .B(KEYINPUT64), .Z(n446) );
  XNOR2_X1 U503 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n456) );
  XOR2_X1 U505 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U508 ( .A(n452), .B(n451), .Z(n454) );
  XNOR2_X1 U509 ( .A(G113GAT), .B(G197GAT), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n458) );
  XOR2_X1 U512 ( .A(n458), .B(n457), .Z(n584) );
  INV_X1 U513 ( .A(n584), .ZN(n553) );
  XOR2_X1 U514 ( .A(KEYINPUT67), .B(n553), .Z(n538) );
  OR2_X1 U515 ( .A1(n465), .A2(n538), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT71), .ZN(n491) );
  NAND2_X1 U517 ( .A1(n521), .A2(n491), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT38), .B(KEYINPUT108), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n461), .B(n460), .ZN(n506) );
  NOR2_X1 U520 ( .A1(n528), .A2(n506), .ZN(n464) );
  INV_X1 U521 ( .A(G218GAT), .ZN(n486) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT41), .ZN(n557) );
  INV_X1 U523 ( .A(n557), .ZN(n540) );
  NAND2_X1 U524 ( .A1(n540), .A2(n584), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n592), .A2(n468), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT118), .ZN(n470) );
  AND2_X1 U527 ( .A1(n470), .A2(n563), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT47), .ZN(n476) );
  NOR2_X1 U529 ( .A1(n483), .A2(n560), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT45), .B(n472), .Z(n473) );
  NOR2_X1 U531 ( .A1(n465), .A2(n473), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n474), .A2(n538), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n533) );
  NOR2_X1 U536 ( .A1(n533), .A2(n524), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT54), .B(n479), .ZN(n569) );
  AND2_X1 U538 ( .A1(n569), .A2(n567), .ZN(n481) );
  INV_X1 U539 ( .A(n480), .ZN(n551) );
  AND2_X1 U540 ( .A1(n481), .A2(n551), .ZN(n593) );
  INV_X1 U541 ( .A(n593), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT62), .B(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1355GAT) );
  NAND2_X1 U545 ( .A1(n592), .A2(n563), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT79), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT16), .ZN(n490) );
  AND2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n510) );
  NAND2_X1 U549 ( .A1(n491), .A2(n510), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n567), .A2(n499), .ZN(n492) );
  XOR2_X1 U551 ( .A(n492), .B(KEYINPUT34), .Z(n493) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n524), .A2(n499), .ZN(n494) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n494), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n499), .A2(n572), .ZN(n498) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n496) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n528), .A2(n499), .ZN(n500) );
  XOR2_X1 U561 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U562 ( .A1(n567), .A2(n506), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n524), .A2(n506), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  NOR2_X1 U569 ( .A1(n572), .A2(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  XNOR2_X1 U573 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n584), .A2(n557), .ZN(n520) );
  AND2_X1 U575 ( .A1(n520), .A2(n510), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT114), .B(n511), .Z(n517) );
  NOR2_X1 U577 ( .A1(n567), .A2(n517), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n517), .A2(n524), .ZN(n515) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n572), .ZN(n516) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  NOR2_X1 U585 ( .A1(n528), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U588 ( .A1(n567), .A2(n527), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n572), .A2(n527), .ZN(n526) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  INV_X1 U599 ( .A(n572), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n552) );
  NAND2_X1 U601 ( .A1(n534), .A2(n552), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT120), .B(n535), .ZN(n536) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n548) );
  INV_X1 U604 ( .A(n538), .ZN(n573) );
  NAND2_X1 U605 ( .A1(n548), .A2(n573), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U608 ( .A1(n548), .A2(n540), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n545) );
  NAND2_X1 U613 ( .A1(n548), .A2(n592), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  INV_X1 U617 ( .A(n563), .ZN(n581) );
  NAND2_X1 U618 ( .A1(n548), .A2(n581), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n553), .A2(n562), .ZN(n554) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n557), .A2(n562), .ZN(n558) );
  XOR2_X1 U627 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  XOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT125), .Z(n575) );
  INV_X1 U633 ( .A(n565), .ZN(n566) );
  AND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  AND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT55), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n575), .B(n574), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n580), .A2(n540), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U643 ( .A1(n580), .A2(n592), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT58), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n588) );
  XOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT126), .Z(n586) );
  NAND2_X1 U650 ( .A1(n593), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U654 ( .A1(n593), .A2(n465), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(G204GAT), .B(n591), .Z(G1353GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
endmodule

