//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G1gat), .B2(new_n207), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(G8gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT87), .B(G43gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  OR2_X1    g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n219), .B2(new_n215), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT88), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n218), .B1(new_n227), .B2(new_n223), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n222), .A2(new_n226), .B1(new_n228), .B2(new_n220), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n220), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n212), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n230), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT13), .Z(new_n239));
  NOR3_X1   g038(.A1(new_n213), .A2(new_n229), .A3(new_n235), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  INV_X1    g042(.A(new_n234), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT89), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n233), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n229), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n212), .B1(new_n233), .B2(new_n246), .ZN(new_n250));
  AOI211_X1 g049(.A(new_n243), .B(new_n244), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n242), .B1(new_n251), .B2(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n238), .A3(new_n234), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n206), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(KEYINPUT18), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  INV_X1    g058(.A(new_n206), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n242), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G155gat), .B(G162gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(KEYINPUT77), .A3(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273));
  INV_X1    g072(.A(new_n269), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n275), .A3(new_n264), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT78), .B(G155gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n268), .B1(new_n277), .B2(G162gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n280));
  AND2_X1   g079(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n282));
  OAI21_X1  g081(.A(G162gat), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n284), .A2(new_n264), .A3(new_n272), .A4(new_n275), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n271), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT1), .ZN(new_n289));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(KEYINPUT1), .B2(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n280), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n279), .B2(new_n294), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n291), .A2(new_n293), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT4), .A3(new_n271), .A4(new_n285), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n295), .A2(new_n296), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n296), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n279), .A2(new_n294), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n285), .A2(new_n271), .B1(new_n291), .B2(new_n293), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n300), .A2(new_n298), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(KEYINPUT5), .A3(new_n296), .A4(new_n295), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT85), .ZN(new_n311));
  XOR2_X1   g110(.A(G1gat), .B(G29gat), .Z(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(new_n309), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n311), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT6), .B1(new_n310), .B2(new_n316), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT6), .A4(new_n317), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  INV_X1    g126(.A(G211gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n326), .A3(new_n330), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  OR2_X1    g137(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT28), .A3(new_n344), .ZN(new_n349));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT26), .ZN(new_n351));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n351), .A2(new_n356), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n347), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359));
  NAND3_X1  g158(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(G183gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n339), .A2(new_n361), .A3(new_n340), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n360), .B(new_n362), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n368), .A2(new_n369), .B1(KEYINPUT23), .B2(new_n350), .ZN(new_n370));
  INV_X1    g169(.A(G169gat), .ZN(new_n371));
  INV_X1    g170(.A(G176gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT25), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n360), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  INV_X1    g177(.A(new_n363), .ZN(new_n379));
  OR2_X1    g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(KEYINPUT65), .A3(new_n360), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n372), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT23), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n354), .A2(new_n355), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(KEYINPUT23), .A3(new_n372), .A4(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n378), .A2(new_n381), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389));
  AOI221_X4 g188(.A(new_n359), .B1(new_n367), .B2(new_n375), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n375), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT70), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n358), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n398), .B(new_n358), .C1(new_n390), .C2(new_n393), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n358), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n405), .B2(new_n396), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n395), .A2(new_n401), .A3(new_n397), .A4(new_n399), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n337), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n397), .A2(KEYINPUT29), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n399), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n358), .A2(new_n397), .A3(new_n402), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n411), .A2(new_n337), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n409), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n325), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n409), .B2(new_n413), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(KEYINPUT37), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n336), .B1(new_n407), .B2(new_n408), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n411), .A2(new_n336), .A3(new_n412), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n408), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n413), .B1(new_n431), .B2(new_n336), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n433), .A2(KEYINPUT37), .B1(new_n421), .B2(new_n422), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n420), .B(new_n430), .C1(new_n434), .C2(new_n424), .ZN(new_n435));
  INV_X1    g234(.A(G22gat), .ZN(new_n436));
  INV_X1    g235(.A(G228gat), .ZN(new_n437));
  INV_X1    g236(.A(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n286), .B1(new_n337), .B2(KEYINPUT29), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n279), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n336), .B1(new_n287), .B2(new_n404), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n279), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n335), .A2(KEYINPUT80), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n404), .C1(new_n336), .C2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n445), .B1(new_n448), .B2(new_n286), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n449), .A2(new_n441), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n436), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n436), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT82), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT31), .B(G50gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n452), .A2(new_n457), .A3(new_n453), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n452), .A2(KEYINPUT83), .A3(new_n457), .A4(new_n453), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n431), .A2(new_n336), .ZN(new_n467));
  INV_X1    g266(.A(new_n413), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n468), .A4(new_n416), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n469), .B(new_n421), .C1(new_n418), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n295), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n300), .A2(new_n298), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n302), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n303), .A2(new_n304), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n475), .B(KEYINPUT39), .C1(new_n302), .C2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n316), .B1(new_n475), .B2(KEYINPUT39), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT40), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n320), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n478), .B(KEYINPUT84), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT40), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n466), .B1(new_n472), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n435), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n322), .B1(new_n316), .B2(new_n310), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n324), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n466), .B1(new_n472), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n394), .A2(new_n294), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n299), .B(new_n358), .C1(new_n390), .C2(new_n393), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT64), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(new_n495), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT34), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT73), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n496), .A2(KEYINPUT34), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n492), .A2(new_n493), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  XOR2_X1   g304(.A(G15gat), .B(G43gat), .Z(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n497), .B2(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n508), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n500), .A2(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n498), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n511), .B1(new_n504), .B2(new_n505), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n517), .A3(new_n514), .ZN(new_n521));
  INV_X1    g320(.A(new_n498), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(KEYINPUT36), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n520), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n487), .A2(new_n491), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n465), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n471), .B1(new_n432), .B2(new_n416), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n489), .A3(new_n421), .A4(new_n469), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT35), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n523), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n325), .A2(new_n419), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n537));
  INV_X1    g336(.A(new_n472), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .A4(new_n465), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n263), .B1(new_n529), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G155gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  XOR2_X1   g344(.A(G57gat), .B(G64gat), .Z(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  INV_X1    g346(.A(G71gat), .ZN(new_n548));
  INV_X1    g347(.A(G78gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(KEYINPUT91), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n212), .B1(KEYINPUT21), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n553), .A2(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G127gat), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n555), .A3(new_n561), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n545), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n560), .A2(new_n561), .A3(new_n555), .ZN(new_n566));
  INV_X1    g365(.A(new_n545), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n566), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT94), .B(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G99gat), .ZN(new_n576));
  INV_X1    g375(.A(G106gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT8), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n579), .A2(new_n581), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT41), .ZN(new_n585));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT92), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n584), .A2(new_n229), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n246), .B2(new_n233), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n249), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT95), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OR3_X1    g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n592), .B1(new_n591), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n587), .A2(new_n585), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n591), .A2(new_n595), .B1(KEYINPUT97), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n596), .A2(new_n605), .A3(new_n597), .A4(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n569), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n580), .A2(KEYINPUT98), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n553), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n553), .A2(new_n609), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n583), .B2(new_n582), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n553), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n612), .ZN(new_n619));
  INV_X1    g418(.A(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n621), .A3(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n608), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n541), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n490), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT99), .B(G1gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1324gat));
  AND2_X1   g433(.A1(new_n541), .A2(new_n472), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G8gat), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n630), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n638), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n643));
  OAI221_X1 g442(.A(new_n637), .B1(new_n638), .B2(new_n640), .C1(new_n642), .C2(new_n643), .ZN(G1325gat));
  AND2_X1   g443(.A1(new_n541), .A2(new_n535), .ZN(new_n645));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n630), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n528), .A2(new_n524), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(new_n646), .ZN(G1326gat));
  AND3_X1   g450(.A1(new_n541), .A2(new_n466), .A3(new_n630), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT101), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NOR2_X1   g454(.A1(new_n530), .A2(new_n472), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n469), .A2(new_n421), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(new_n531), .A3(new_n490), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n535), .A2(new_n658), .A3(new_n465), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n656), .A2(new_n537), .B1(new_n659), .B2(KEYINPUT35), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT37), .B1(new_n409), .B2(new_n413), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n424), .B1(new_n423), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n428), .B1(new_n421), .B2(new_n422), .ZN(new_n663));
  INV_X1    g462(.A(new_n419), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n467), .A2(new_n468), .A3(new_n416), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n324), .A4(new_n323), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n485), .B1(new_n657), .B2(new_n531), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n465), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n528), .A2(new_n491), .A3(new_n524), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT102), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n648), .A2(new_n673), .A3(new_n487), .A4(new_n491), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n660), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n607), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n607), .B1(new_n529), .B2(new_n540), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n675), .A2(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n569), .A2(new_n629), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n262), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n489), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n682), .A2(G29gat), .A3(new_n489), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(G1328gat));
  INV_X1    g488(.A(G36gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n681), .A2(new_n676), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n635), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT46), .Z(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n684), .B2(new_n538), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1329gat));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n672), .A2(new_n674), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n678), .B1(new_n698), .B2(new_n540), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n677), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n649), .B(new_n683), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n216), .ZN(new_n702));
  INV_X1    g501(.A(new_n216), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n645), .A2(new_n703), .A3(new_n692), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n697), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n697), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT103), .B(new_n708), .C1(new_n702), .C2(new_n704), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n680), .A2(new_n466), .A3(new_n683), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n680), .A2(KEYINPUT106), .A3(new_n466), .A4(new_n683), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(G50gat), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n691), .A2(G50gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n541), .A2(new_n466), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT48), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n711), .A2(G50gat), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n717), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n715), .A2(new_n719), .B1(new_n721), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g521(.A1(new_n565), .A2(new_n568), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n676), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n263), .A3(new_n629), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n675), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n490), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g527(.A1(new_n675), .A2(new_n538), .A3(new_n725), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  AOI21_X1  g532(.A(new_n548), .B1(new_n726), .B2(new_n649), .ZN(new_n734));
  AOI21_X1  g533(.A(G71gat), .B1(new_n519), .B2(new_n523), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g536(.A1(new_n726), .A2(new_n466), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(new_n629), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n569), .A2(new_n262), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n680), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n489), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT102), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n528), .A2(new_n491), .A3(new_n524), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n673), .B1(new_n745), .B2(new_n487), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n540), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n569), .A2(new_n262), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n676), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n675), .B2(new_n749), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n490), .A2(new_n574), .A3(new_n629), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT107), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n743), .B1(new_n756), .B2(new_n758), .ZN(G1336gat));
  AND3_X1   g558(.A1(new_n680), .A2(new_n472), .A3(new_n741), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n538), .A2(G92gat), .A3(new_n740), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n751), .B2(new_n754), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n760), .A2(new_n573), .B1(new_n763), .B2(KEYINPUT108), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(new_n573), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n742), .B2(new_n538), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n767), .A2(new_n768), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n742), .B2(new_n648), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n535), .A2(new_n576), .A3(new_n629), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n756), .B2(new_n775), .ZN(G1338gat));
  OAI21_X1  g575(.A(G106gat), .B1(new_n742), .B2(new_n465), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n465), .A2(G106gat), .A3(new_n740), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n752), .B2(new_n755), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT53), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n777), .B(new_n779), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1339gat));
  AOI21_X1  g585(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n787), .B2(new_n238), .ZN(new_n788));
  INV_X1    g587(.A(new_n239), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n236), .B2(new_n240), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n787), .A2(KEYINPUT112), .A3(new_n238), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n205), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n261), .A3(new_n629), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n614), .A2(new_n620), .A3(new_n615), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n618), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n620), .B1(new_n614), .B2(new_n615), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n625), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n628), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n262), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g605(.A(KEYINPUT111), .B(KEYINPUT55), .C1(new_n796), .C2(new_n799), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n794), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n607), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n801), .A2(new_n604), .A3(new_n606), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n261), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n811), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n569), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n569), .A2(new_n263), .A3(new_n607), .A4(new_n740), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n262), .B(new_n801), .C1(new_n806), .C2(new_n807), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n676), .B1(new_n818), .B2(new_n794), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n811), .A2(new_n808), .A3(new_n812), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n723), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(new_n815), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n489), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n656), .ZN(new_n826));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n262), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n824), .A2(new_n466), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n538), .A2(new_n490), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n535), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(G113gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n832), .A3(new_n263), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n833), .ZN(G1340gat));
  AOI21_X1  g633(.A(G120gat), .B1(new_n826), .B2(new_n629), .ZN(new_n835));
  INV_X1    g634(.A(G120gat), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n831), .A2(new_n836), .A3(new_n740), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(G1341gat));
  NAND3_X1  g637(.A1(new_n826), .A2(new_n559), .A3(new_n569), .ZN(new_n839));
  OAI21_X1  g638(.A(G127gat), .B1(new_n831), .B2(new_n723), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n607), .A2(G134gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n831), .B2(new_n607), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n825), .A2(new_n656), .ZN(new_n846));
  INV_X1    g645(.A(new_n843), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT56), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n844), .A2(new_n845), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1343gat));
  AND2_X1   g652(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n648), .A2(new_n466), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n472), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(new_n817), .A3(new_n490), .A4(new_n823), .ZN(new_n857));
  INV_X1    g656(.A(G141gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n262), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT118), .Z(new_n860));
  NOR2_X1   g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n649), .A2(new_n829), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n824), .B2(new_n465), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n794), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n804), .A2(new_n805), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n262), .A2(new_n801), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n793), .A2(KEYINPUT115), .A3(new_n629), .A4(new_n261), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n607), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n569), .B1(new_n874), .B2(new_n813), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n815), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT57), .B(new_n466), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n865), .B1(new_n867), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n262), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n863), .B1(new_n881), .B2(new_n858), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n861), .A2(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n857), .B2(new_n860), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n858), .B1(new_n880), .B2(new_n262), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(KEYINPUT117), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n882), .B1(new_n888), .B2(new_n862), .ZN(G1344gat));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n629), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n466), .A4(new_n823), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n724), .A2(KEYINPUT120), .A3(new_n263), .A4(new_n740), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n815), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n466), .B1(new_n875), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n866), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT59), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT121), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n902), .B(KEYINPUT59), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n880), .A2(new_n629), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n857), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n899), .A3(new_n629), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1345gat));
  AOI21_X1  g710(.A(new_n277), .B1(new_n909), .B2(new_n569), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n569), .A2(new_n277), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT122), .Z(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n880), .B2(new_n914), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n909), .B2(new_n676), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n676), .A2(G162gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n880), .B2(new_n917), .ZN(G1347gat));
  NAND4_X1  g717(.A1(new_n828), .A2(new_n489), .A3(new_n472), .A4(new_n535), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n263), .ZN(new_n920));
  NOR4_X1   g719(.A1(new_n824), .A2(new_n490), .A3(new_n538), .A4(new_n530), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(new_n385), .A3(new_n386), .A4(new_n262), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n919), .B2(new_n740), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n372), .A3(new_n629), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n919), .B2(new_n723), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n343), .A3(new_n569), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n921), .A2(new_n341), .A3(new_n676), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n919), .A2(new_n607), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(G190gat), .ZN(new_n938));
  OAI211_X1 g737(.A(G190gat), .B(new_n936), .C1(new_n919), .C2(new_n607), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n938), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n855), .A2(new_n538), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n942), .A2(new_n817), .A3(new_n489), .A4(new_n823), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n262), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n648), .A2(new_n489), .A3(new_n472), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n891), .B2(new_n897), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n262), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(new_n947), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n950), .B2(new_n740), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n740), .A2(G204gat), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n943), .A2(KEYINPUT62), .A3(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n328), .A3(new_n569), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n723), .B(new_n946), .C1(new_n891), .C2(new_n897), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n328), .B1(new_n957), .B2(KEYINPUT125), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT125), .B1(new_n947), .B2(new_n569), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n891), .A2(new_n897), .ZN(new_n962));
  INV_X1    g761(.A(new_n946), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n569), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G211gat), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(new_n959), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n956), .B1(new_n961), .B2(new_n967), .ZN(G1354gat));
  OAI21_X1  g767(.A(new_n329), .B1(new_n943), .B2(new_n607), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n607), .A2(new_n329), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n950), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


