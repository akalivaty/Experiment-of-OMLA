//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G2106), .B2(new_n453), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(new_n468), .B2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n461), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT66), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n469), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n479), .A2(new_n469), .A3(new_n480), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n480), .B1(new_n479), .B2(new_n469), .ZN(new_n489));
  OAI21_X1  g064(.A(G125), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n483), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n474), .B1(new_n487), .B2(new_n492), .ZN(G160));
  NAND4_X1  g068(.A1(new_n471), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n461), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G136), .ZN(new_n499));
  OAI221_X1 g074(.A(new_n496), .B1(new_n497), .B2(new_n498), .C1(new_n499), .C2(new_n472), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT71), .A2(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT71), .A2(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n461), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n494), .A2(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n471), .A2(new_n467), .A3(new_n469), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n508), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n488), .B2(new_n489), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n507), .B1(new_n511), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(G62), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n518), .A2(new_n519), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n515), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT6), .A3(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n523), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G50), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n524), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n528), .A2(new_n539), .ZN(G166));
  NAND3_X1  g115(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n533), .A2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n541), .B(new_n542), .C1(new_n546), .C2(KEYINPUT74), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(G168));
  AOI22_X1  g124(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n516), .A2(new_n517), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n530), .B2(new_n532), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G90), .B1(G52), .B2(new_n533), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(G171));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n555), .A2(G81), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n533), .A2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n538), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G91), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n533), .A2(new_n575), .A3(G53), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n537), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n515), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n577), .A3(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n573), .A2(G87), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n537), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G49), .B2(new_n533), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n554), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n533), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n555), .A2(new_n572), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n554), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n555), .A2(G85), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n533), .A2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  INV_X1    g179(.A(new_n533), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(new_n605), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(G66), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(G66), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n537), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n523), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT10), .B1(new_n573), .B2(G92), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n573), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(G868), .B2(new_n624), .ZN(G297));
  XOR2_X1   g200(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n478), .A2(new_n481), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n463), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n640), .A2(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(new_n640), .ZN(new_n644));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n494), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G135), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(new_n472), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n638), .A2(new_n639), .A3(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1341), .B(G1348), .Z(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  AOI21_X1  g250(.A(KEYINPUT18), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(new_n677));
  NOR2_X1   g252(.A1(G2072), .A2(G2078), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n442), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n673), .B2(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2096), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT87), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT87), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n687), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n693), .C1(new_n685), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(KEYINPUT97), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n566), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n704), .B2(G19), .ZN(new_n706));
  INV_X1    g281(.A(G1341), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G171), .A2(new_n704), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G5), .B2(new_n704), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G33), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  INV_X1    g290(.A(G139), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n472), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n633), .A2(G127), .ZN(new_n718));
  INV_X1    g293(.A(G115), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n466), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(new_n712), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n710), .A2(new_n711), .B1(G2072), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n706), .A2(new_n707), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G28), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n712), .B1(new_n725), .B2(G28), .ZN(new_n727));
  AND2_X1   g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NOR2_X1   g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n649), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G29), .ZN(new_n732));
  AND4_X1   g307(.A1(new_n708), .A2(new_n723), .A3(new_n724), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n710), .A2(new_n711), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n704), .A2(G20), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT23), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n624), .B2(new_n704), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G1956), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n704), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n704), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n712), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n495), .A2(G129), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n463), .A2(G105), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n472), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(G141), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(new_n712), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n722), .A2(G2072), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n733), .A2(new_n741), .A3(new_n745), .A4(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n734), .A2(new_n735), .B1(G1956), .B2(new_n739), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT91), .ZN(new_n763));
  INV_X1    g338(.A(new_n619), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n608), .B(new_n615), .C1(new_n764), .C2(new_n617), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n763), .B1(new_n765), .B2(new_n704), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1348), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n712), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n712), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G2078), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n712), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n774));
  INV_X1    g349(.A(G128), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n494), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n752), .B2(G140), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(new_n712), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n761), .A2(new_n767), .A3(new_n770), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n760), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g358(.A1(G162), .A2(G29), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G29), .B2(G35), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n783), .B(new_n791), .C1(new_n788), .C2(new_n789), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n782), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n790), .A2(new_n791), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n712), .B1(KEYINPUT24), .B2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(KEYINPUT24), .B2(G34), .ZN(new_n798));
  INV_X1    g373(.A(G160), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT92), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n796), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n703), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n794), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n792), .A2(new_n760), .A3(new_n808), .A4(new_n781), .ZN(new_n809));
  INV_X1    g384(.A(new_n806), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT97), .ZN(new_n811));
  NOR2_X1   g386(.A1(G25), .A2(G29), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n814));
  INV_X1    g389(.A(G119), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n494), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n752), .B2(G131), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n812), .B1(new_n817), .B2(G29), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  OAI21_X1  g395(.A(KEYINPUT90), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n704), .A2(G24), .ZN(new_n822));
  INV_X1    g397(.A(G290), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n704), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G1986), .Z(new_n826));
  AOI211_X1 g401(.A(new_n821), .B(new_n826), .C1(new_n819), .C2(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n704), .A2(G23), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n584), .A2(new_n586), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n704), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT33), .ZN(new_n831));
  INV_X1    g406(.A(G1976), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  MUX2_X1   g408(.A(G6), .B(G305), .S(G16), .Z(new_n834));
  XOR2_X1   g409(.A(KEYINPUT32), .B(G1981), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G22), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n837), .A2(KEYINPUT89), .A3(G16), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT89), .B1(new_n837), .B2(G16), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n838), .B(new_n839), .C1(G166), .C2(new_n704), .ZN(new_n840));
  INV_X1    g415(.A(G1971), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n833), .A2(KEYINPUT34), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT34), .B1(new_n833), .B2(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n827), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n827), .A2(new_n844), .A3(new_n848), .A4(new_n845), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n807), .A2(new_n811), .B1(new_n847), .B2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n807), .A2(new_n811), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(G150));
  AOI22_X1  g428(.A1(new_n555), .A2(G93), .B1(G55), .B2(new_n533), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT98), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n515), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NOR2_X1   g435(.A1(new_n765), .A2(new_n627), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n566), .A3(new_n857), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n566), .B1(new_n855), .B2(new_n857), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n753), .B(new_n721), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n495), .A2(G130), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n461), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(G142), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n876), .B1(new_n877), .B2(new_n878), .C1(new_n879), .C2(new_n472), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n635), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n875), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n777), .B(G164), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n817), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n884), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(new_n731), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G160), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n886), .A2(new_n887), .B1(new_n889), .B2(KEYINPUT101), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(KEYINPUT101), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n882), .A2(new_n884), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n885), .ZN(new_n894));
  INV_X1    g469(.A(new_n889), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT100), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(KEYINPUT100), .A3(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g474(.A1(new_n765), .A2(new_n624), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n620), .A2(G299), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n620), .A2(G299), .A3(KEYINPUT102), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n866), .B(new_n629), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  XNOR2_X1  g488(.A(G288), .B(G166), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n823), .B(G305), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n914), .B(new_n915), .Z(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n910), .B(new_n918), .C1(new_n909), .C2(new_n911), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n913), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n858), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(G868), .B2(new_n923), .ZN(G295));
  OAI21_X1  g499(.A(new_n922), .B1(G868), .B2(new_n923), .ZN(G331));
  AOI21_X1  g500(.A(G171), .B1(G286), .B2(KEYINPUT104), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n858), .A2(new_n565), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g504(.A1(G168), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n930), .A3(new_n863), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n928), .B2(new_n863), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n929), .B(G168), .C1(new_n864), .C2(new_n865), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n926), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n908), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n911), .B2(new_n937), .ZN(new_n939));
  INV_X1    g514(.A(new_n916), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n938), .B(new_n916), .C1(new_n911), .C2(new_n937), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n900), .A2(new_n901), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n906), .B1(new_n934), .B2(new_n936), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n945), .B(new_n916), .C1(new_n911), .C2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n937), .A2(new_n911), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n936), .A2(new_n934), .B1(new_n905), .B2(new_n907), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n940), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g526(.A1(KEYINPUT43), .A2(new_n947), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT44), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n955), .A2(new_n947), .A3(new_n948), .A4(new_n951), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(G397));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n963), .B(new_n474), .C1(new_n487), .C2(new_n492), .ZN(new_n964));
  INV_X1    g539(.A(new_n507), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n513), .A2(new_n511), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(KEYINPUT105), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n969), .B2(KEYINPUT105), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n962), .B1(new_n972), .B2(G1996), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n972), .A2(new_n962), .A3(G1996), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n961), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n975), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(KEYINPUT46), .A3(new_n973), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT125), .ZN(new_n980));
  INV_X1    g555(.A(new_n972), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n777), .B(G2067), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n753), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n980), .B1(new_n979), .B2(new_n984), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n960), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n987), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT47), .A3(new_n985), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n753), .B1(new_n974), .B2(new_n975), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n982), .B1(new_n992), .B2(new_n753), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n981), .A2(new_n993), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n817), .A2(new_n991), .A3(new_n820), .A4(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n777), .A2(new_n779), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n981), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n817), .B(new_n820), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n981), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT126), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G290), .A2(G1986), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT106), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n981), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1009));
  AND4_X1   g584(.A1(new_n988), .A2(new_n990), .A3(new_n997), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n633), .A2(new_n512), .B1(KEYINPUT4), .B2(new_n510), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT45), .B(new_n968), .C1(new_n1014), .C2(new_n507), .ZN(new_n1015));
  NAND4_X1  g590(.A1(G160), .A2(G40), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1011), .B1(new_n1016), .B2(G2078), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n968), .C1(new_n1014), .C2(new_n507), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n487), .A2(new_n492), .ZN(new_n1024));
  INV_X1    g599(.A(new_n474), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1023), .A2(new_n1024), .A3(G40), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n711), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1021), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n967), .B2(new_n968), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1012), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1011), .A2(G2078), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n964), .A3(new_n1015), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1017), .A2(new_n1027), .A3(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1033), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT123), .B1(new_n1033), .B2(G171), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT55), .B(G8), .C1(new_n528), .C2(new_n539), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT110), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  INV_X1    g614(.A(new_n527), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G75), .A2(G543), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n526), .B2(KEYINPUT73), .ZN(new_n1042));
  OAI21_X1  g617(.A(G651), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n555), .A2(G88), .B1(G50), .B2(new_n533), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT111), .B1(new_n1045), .B2(KEYINPUT55), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1047), .B(new_n1048), .C1(G166), .C2(new_n1039), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1019), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1019), .B(new_n968), .C1(new_n1014), .C2(new_n507), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1024), .A2(G40), .A3(new_n1025), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1055), .A2(new_n791), .B1(new_n841), .B2(new_n1016), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1051), .B1(new_n1056), .B2(new_n1039), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n591), .B1(new_n595), .B2(new_n538), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G1981), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1061), .A3(KEYINPUT49), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT49), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(G160), .A2(G40), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(G8), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n584), .A2(G1976), .A3(new_n586), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(G288), .B2(new_n832), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1065), .A2(G8), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT67), .B1(new_n491), .B2(G2105), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n486), .B(new_n461), .C1(new_n490), .C2(new_n483), .ZN(new_n1072));
  OAI211_X1 g647(.A(G40), .B(new_n1025), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1067), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1066), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1016), .A2(new_n841), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n964), .A2(new_n1078), .A3(new_n791), .A4(new_n1023), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1037), .B(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1039), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1080), .A2(new_n1084), .A3(KEYINPUT112), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT112), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1057), .B(new_n1076), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1036), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT45), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1024), .A2(G40), .A3(new_n1025), .A4(new_n1015), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n744), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n964), .A2(new_n1078), .A3(new_n801), .A4(new_n1023), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(G168), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT62), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1101), .A3(new_n1098), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1088), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1076), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1080), .A2(new_n1084), .A3(KEYINPUT112), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1039), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1053), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1073), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT50), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n791), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1039), .B1(new_n1115), .B2(new_n1077), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1051), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1110), .B(new_n1111), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1104), .B1(new_n1109), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1051), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1110), .A2(new_n1121), .A3(G168), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1122), .B2(new_n1076), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n829), .A2(new_n832), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT113), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1039), .B(new_n1124), .C1(new_n1127), .C2(new_n1059), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1119), .A2(new_n1123), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1103), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1133));
  OR2_X1    g708(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n964), .A2(new_n1013), .A3(new_n1015), .A4(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1348), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1124), .A2(new_n779), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n765), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT114), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1134), .A2(new_n1133), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1956), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1135), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1016), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1137), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1148), .B2(new_n1137), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1148), .B2(new_n1137), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  OAI22_X1  g730(.A1(KEYINPUT120), .A2(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1148), .A2(new_n1137), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1153), .B(KEYINPUT61), .C1(new_n1157), .C2(new_n1151), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n620), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1139), .A2(new_n1161), .A3(new_n1140), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n620), .A2(new_n1160), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT60), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1162), .B1(new_n1165), .B2(new_n1163), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1164), .A2(new_n1166), .A3(KEYINPUT122), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT122), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1156), .B(new_n1158), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT115), .B(G1996), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n964), .A2(new_n1013), .A3(new_n1015), .A4(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT58), .B(G1341), .Z(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1172), .A2(KEYINPUT116), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT116), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n566), .B(new_n1170), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1177), .A2(KEYINPUT118), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n566), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1177), .A2(KEYINPUT118), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1150), .B1(new_n1169), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1027), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(KEYINPUT124), .B(new_n711), .C1(new_n1022), .C2(new_n1026), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n970), .A2(new_n971), .ZN(new_n1187));
  AND4_X1   g762(.A1(G40), .A2(new_n1025), .A3(new_n485), .A4(new_n1031), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(new_n1015), .A3(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1185), .A2(new_n1186), .A3(new_n1017), .A4(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1190), .A2(G171), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT54), .B1(new_n1036), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT54), .B1(new_n1033), .B2(G171), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1194), .B1(G171), .B2(new_n1190), .ZN(new_n1195));
  NOR4_X1   g770(.A1(new_n1192), .A2(new_n1193), .A3(new_n1087), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1130), .B1(new_n1183), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1006), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT107), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1200), .A2(new_n1000), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1010), .B1(new_n1197), .B2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g777(.A1(new_n668), .A2(G319), .ZN(new_n1204));
  NOR3_X1   g778(.A1(G229), .A2(G227), .A3(new_n1204), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n1205), .B(new_n898), .C1(new_n956), .C2(new_n957), .ZN(G225));
  INV_X1    g780(.A(G225), .ZN(G308));
endmodule


