// Benchmark "locked_c1908" written by ABC on Sat Dec 16 10:46:12 2023

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n441, new_n442, new_n443, new_n444, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n485,
    new_n486, new_n487, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n520,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n123));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n124));
  XNOR2_X1  g002(.A(new_n123), .B(new_n124), .ZN(new_n125));
  INV_X1    g003(.A(new_n125), .ZN(new_n126));
  INV_X1    g004(.A(G131), .ZN(new_n127));
  INV_X1    g005(.A(G137), .ZN(new_n128));
  NAND3_X1  g006(.A1(new_n128), .A2(KEYINPUT11), .A3(G134), .ZN(new_n129));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n130));
  INV_X1    g008(.A(G134), .ZN(new_n131));
  AOI21_X1  g009(.A(new_n130), .B1(new_n131), .B2(G137), .ZN(new_n132));
  NOR2_X1   g010(.A1(new_n131), .A2(G137), .ZN(new_n133));
  OAI211_X1 g011(.A(new_n127), .B(new_n129), .C1(new_n132), .C2(new_n133), .ZN(new_n134));
  INV_X1    g012(.A(G143), .ZN(new_n135));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n135), .B2(G146), .ZN(new_n136));
  NOR2_X1   g014(.A1(new_n135), .A2(G146), .ZN(new_n137));
  INV_X1    g015(.A(G146), .ZN(new_n138));
  NOR2_X1   g016(.A1(new_n138), .A2(G143), .ZN(new_n139));
  OAI211_X1 g017(.A(G128), .B(new_n136), .C1(new_n137), .C2(new_n139), .ZN(new_n140));
  NAND2_X1  g018(.A1(new_n138), .A2(G143), .ZN(new_n141));
  NAND2_X1  g019(.A1(new_n135), .A2(G146), .ZN(new_n142));
  INV_X1    g020(.A(G128), .ZN(new_n143));
  OAI211_X1 g021(.A(new_n141), .B(new_n142), .C1(KEYINPUT1), .C2(new_n143), .ZN(new_n144));
  NOR2_X1   g022(.A1(new_n128), .A2(G134), .ZN(new_n145));
  OAI21_X1  g023(.A(G131), .B1(new_n133), .B2(new_n145), .ZN(new_n146));
  NAND4_X1  g024(.A1(new_n134), .A2(new_n140), .A3(new_n144), .A4(new_n146), .ZN(new_n147));
  INV_X1    g025(.A(new_n134), .ZN(new_n148));
  OAI21_X1  g026(.A(KEYINPUT11), .B1(new_n128), .B2(G134), .ZN(new_n149));
  NAND2_X1  g027(.A1(new_n128), .A2(G134), .ZN(new_n150));
  NAND2_X1  g028(.A1(new_n149), .A2(new_n150), .ZN(new_n151));
  AOI21_X1  g029(.A(new_n127), .B1(new_n151), .B2(new_n129), .ZN(new_n152));
  NOR2_X1   g030(.A1(new_n148), .A2(new_n152), .ZN(new_n153));
  INV_X1    g031(.A(KEYINPUT0), .ZN(new_n154));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n155));
  OAI21_X1  g033(.A(new_n154), .B1(new_n155), .B2(new_n143), .ZN(new_n156));
  NAND2_X1  g034(.A1(new_n155), .A2(new_n143), .ZN(new_n157));
  OAI211_X1 g035(.A(KEYINPUT0), .B(G128), .C1(new_n137), .C2(new_n139), .ZN(new_n158));
  AND3_X1   g036(.A1(new_n156), .A2(new_n157), .A3(new_n158), .ZN(new_n159));
  OAI21_X1  g037(.A(new_n147), .B1(new_n153), .B2(new_n159), .ZN(new_n160));
  NAND2_X1  g038(.A1(new_n160), .A2(KEYINPUT30), .ZN(new_n161));
  NAND3_X1  g039(.A1(new_n156), .A2(new_n157), .A3(new_n158), .ZN(new_n162));
  OAI21_X1  g040(.A(new_n162), .B1(new_n148), .B2(new_n152), .ZN(new_n163));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n164));
  NAND3_X1  g042(.A1(new_n163), .A2(new_n164), .A3(new_n147), .ZN(new_n165));
  AOI21_X1  g043(.A(new_n126), .B1(new_n161), .B2(new_n165), .ZN(new_n166));
  NAND3_X1  g044(.A1(new_n163), .A2(new_n126), .A3(new_n147), .ZN(new_n167));
  NOR2_X1   g045(.A1(G237), .A2(G953), .ZN(new_n168));
  NAND2_X1  g046(.A1(new_n168), .A2(G210), .ZN(new_n169));
  XNOR2_X1  g047(.A(new_n169), .B(KEYINPUT27), .ZN(new_n170));
  XNOR2_X1  g048(.A(KEYINPUT26), .B(G101), .ZN(new_n171));
  XNOR2_X1  g049(.A(new_n170), .B(new_n171), .ZN(new_n172));
  NAND2_X1  g050(.A1(new_n167), .A2(new_n172), .ZN(new_n173));
  OAI21_X1  g051(.A(KEYINPUT31), .B1(new_n166), .B2(new_n173), .ZN(new_n174));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n175));
  NAND2_X1  g053(.A1(new_n167), .A2(new_n175), .ZN(new_n176));
  NAND2_X1  g054(.A1(new_n160), .A2(new_n125), .ZN(new_n177));
  NAND4_X1  g055(.A1(new_n163), .A2(new_n126), .A3(KEYINPUT28), .A4(new_n147), .ZN(new_n178));
  NAND3_X1  g056(.A1(new_n176), .A2(new_n177), .A3(new_n178), .ZN(new_n179));
  INV_X1    g057(.A(new_n172), .ZN(new_n180));
  NAND2_X1  g058(.A1(new_n179), .A2(new_n180), .ZN(new_n181));
  AND3_X1   g059(.A1(new_n163), .A2(new_n164), .A3(new_n147), .ZN(new_n182));
  AOI21_X1  g060(.A(new_n164), .B1(new_n163), .B2(new_n147), .ZN(new_n183));
  OAI21_X1  g061(.A(new_n125), .B1(new_n182), .B2(new_n183), .ZN(new_n184));
  INV_X1    g062(.A(KEYINPUT31), .ZN(new_n185));
  INV_X1    g063(.A(new_n173), .ZN(new_n186));
  NAND3_X1  g064(.A1(new_n184), .A2(new_n185), .A3(new_n186), .ZN(new_n187));
  NAND3_X1  g065(.A1(new_n174), .A2(new_n181), .A3(new_n187), .ZN(new_n188));
  NOR2_X1   g066(.A1(G472), .A2(G902), .ZN(new_n189));
  NAND2_X1  g067(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n191));
  NAND2_X1  g069(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  AOI21_X1  g070(.A(new_n172), .B1(new_n184), .B2(new_n167), .ZN(new_n193));
  NAND4_X1  g071(.A1(new_n176), .A2(new_n177), .A3(new_n172), .A4(new_n178), .ZN(new_n194));
  INV_X1    g072(.A(new_n194), .ZN(new_n195));
  NOR3_X1   g073(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT29), .ZN(new_n196));
  INV_X1    g074(.A(G902), .ZN(new_n197));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n198));
  OAI21_X1  g076(.A(new_n197), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g077(.A(G472), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g078(.A1(new_n188), .A2(KEYINPUT32), .A3(new_n189), .ZN(new_n201));
  NAND3_X1  g079(.A1(new_n192), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g081(.A(G119), .ZN(new_n204));
  OAI21_X1  g082(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND3_X1  g083(.A1(new_n143), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  OAI211_X1 g084(.A(new_n205), .B(new_n206), .C1(G119), .C2(new_n143), .ZN(new_n207));
  NAND2_X1  g085(.A1(new_n207), .A2(G110), .ZN(new_n208));
  XOR2_X1   g086(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  XNOR2_X1  g087(.A(G119), .B(G128), .ZN(new_n210));
  NAND2_X1  g088(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g089(.A(G125), .B(G140), .ZN(new_n212));
  NAND2_X1  g090(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n213));
  INV_X1    g091(.A(G140), .ZN(new_n214));
  NAND2_X1  g092(.A1(new_n214), .A2(G125), .ZN(new_n215));
  OR2_X1    g093(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  AND3_X1   g094(.A1(new_n213), .A2(G146), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g095(.A(G146), .B1(new_n213), .B2(new_n216), .ZN(new_n218));
  OAI211_X1 g096(.A(new_n208), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI22_X1  g097(.A1(new_n207), .A2(G110), .B1(new_n210), .B2(new_n209), .ZN(new_n220));
  NAND3_X1  g098(.A1(new_n213), .A2(G146), .A3(new_n216), .ZN(new_n221));
  INV_X1    g099(.A(G125), .ZN(new_n222));
  NAND2_X1  g100(.A1(new_n222), .A2(G140), .ZN(new_n223));
  NAND2_X1  g101(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g102(.A(new_n220), .B(new_n221), .C1(G146), .C2(new_n224), .ZN(new_n225));
  XOR2_X1   g103(.A(KEYINPUT22), .B(G137), .Z(new_n226));
  INV_X1    g104(.A(G953), .ZN(new_n227));
  NAND3_X1  g105(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g106(.A(new_n226), .B(new_n228), .ZN(new_n229));
  AND3_X1   g107(.A1(new_n219), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g108(.A(new_n229), .B1(new_n219), .B2(new_n225), .ZN(new_n231));
  OAI21_X1  g109(.A(new_n197), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g110(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  INV_X1    g111(.A(G217), .ZN(new_n234));
  AOI21_X1  g112(.A(new_n234), .B1(G234), .B2(new_n197), .ZN(new_n235));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n236));
  OAI211_X1 g114(.A(new_n236), .B(new_n197), .C1(new_n230), .C2(new_n231), .ZN(new_n237));
  NAND3_X1  g115(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  OR2_X1    g116(.A1(new_n230), .A2(new_n231), .ZN(new_n239));
  NOR2_X1   g117(.A1(new_n235), .A2(G902), .ZN(new_n240));
  NAND2_X1  g118(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g119(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g120(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n244));
  OAI21_X1  g122(.A(G221), .B1(new_n244), .B2(G902), .ZN(new_n245));
  INV_X1    g123(.A(new_n245), .ZN(new_n246));
  INV_X1    g124(.A(G101), .ZN(new_n247));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g126(.A(G107), .ZN(new_n249));
  NAND3_X1  g127(.A1(new_n248), .A2(new_n249), .A3(G104), .ZN(new_n250));
  INV_X1    g128(.A(G104), .ZN(new_n251));
  AOI21_X1  g129(.A(KEYINPUT3), .B1(new_n251), .B2(G107), .ZN(new_n252));
  NOR2_X1   g130(.A1(new_n251), .A2(G107), .ZN(new_n253));
  OAI211_X1 g131(.A(new_n247), .B(new_n250), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NOR2_X1   g132(.A1(new_n249), .A2(G104), .ZN(new_n255));
  OAI21_X1  g133(.A(G101), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g134(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g135(.A(new_n257), .ZN(new_n258));
  NAND4_X1  g136(.A1(new_n258), .A2(KEYINPUT10), .A3(new_n144), .A4(new_n140), .ZN(new_n259));
  NAND4_X1  g137(.A1(new_n254), .A2(new_n140), .A3(new_n144), .A4(new_n256), .ZN(new_n260));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n261));
  NAND2_X1  g139(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g140(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n263));
  AND3_X1   g141(.A1(new_n263), .A2(KEYINPUT4), .A3(G101), .ZN(new_n264));
  AOI21_X1  g142(.A(KEYINPUT4), .B1(new_n263), .B2(G101), .ZN(new_n265));
  INV_X1    g143(.A(new_n254), .ZN(new_n266));
  NOR3_X1   g144(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI211_X1 g145(.A(new_n259), .B(new_n262), .C1(new_n267), .C2(new_n159), .ZN(new_n268));
  INV_X1    g146(.A(new_n152), .ZN(new_n269));
  NAND2_X1  g147(.A1(new_n269), .A2(new_n134), .ZN(new_n270));
  NAND2_X1  g148(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g149(.A1(new_n263), .A2(G101), .ZN(new_n272));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n273));
  NAND2_X1  g151(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g152(.A1(new_n263), .A2(KEYINPUT4), .A3(G101), .ZN(new_n275));
  NAND3_X1  g153(.A1(new_n274), .A2(new_n254), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g154(.A1(new_n276), .A2(new_n162), .ZN(new_n277));
  NAND4_X1  g155(.A1(new_n277), .A2(new_n153), .A3(new_n259), .A4(new_n262), .ZN(new_n278));
  XNOR2_X1  g156(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g157(.A(G227), .ZN(new_n280));
  NOR2_X1   g158(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XOR2_X1   g159(.A(new_n279), .B(new_n281), .Z(new_n282));
  AND2_X1   g160(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g161(.A1(new_n140), .A2(new_n144), .ZN(new_n284));
  NAND2_X1  g162(.A1(new_n257), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g163(.A1(new_n285), .A2(new_n260), .ZN(new_n286));
  AOI21_X1  g164(.A(KEYINPUT12), .B1(new_n286), .B2(new_n270), .ZN(new_n287));
  AND3_X1   g165(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n270), .ZN(new_n288));
  OAI21_X1  g166(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g167(.A(new_n282), .ZN(new_n290));
  AOI22_X1  g168(.A1(new_n271), .A2(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g169(.A(G469), .B1(new_n291), .B2(G902), .ZN(new_n292));
  INV_X1    g170(.A(G469), .ZN(new_n293));
  INV_X1    g171(.A(new_n260), .ZN(new_n294));
  AOI22_X1  g172(.A1(new_n254), .A2(new_n256), .B1(new_n140), .B2(new_n144), .ZN(new_n295));
  OAI21_X1  g173(.A(new_n270), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g174(.A(KEYINPUT12), .ZN(new_n297));
  NAND2_X1  g175(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g176(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n270), .ZN(new_n299));
  NAND2_X1  g177(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g178(.A1(new_n300), .A2(new_n278), .A3(new_n282), .ZN(new_n301));
  AOI21_X1  g179(.A(new_n282), .B1(new_n271), .B2(new_n278), .ZN(new_n302));
  OAI211_X1 g180(.A(new_n293), .B(new_n197), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g181(.A(new_n246), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g182(.A1(new_n202), .A2(new_n243), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g183(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g184(.A(new_n306), .ZN(new_n307));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n308));
  INV_X1    g186(.A(G116), .ZN(new_n309));
  OAI21_X1  g187(.A(new_n308), .B1(new_n309), .B2(G119), .ZN(new_n310));
  NAND2_X1  g188(.A1(new_n309), .A2(G119), .ZN(new_n311));
  NAND3_X1  g189(.A1(new_n204), .A2(KEYINPUT5), .A3(G116), .ZN(new_n312));
  NAND3_X1  g190(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g191(.A1(new_n313), .A2(G113), .ZN(new_n314));
  NAND2_X1  g192(.A1(new_n123), .A2(new_n124), .ZN(new_n315));
  NAND2_X1  g193(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI22_X1  g194(.A1(new_n267), .A2(new_n126), .B1(new_n257), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g195(.A(G110), .B(G122), .Z(new_n318));
  NAND3_X1  g196(.A1(new_n317), .A2(KEYINPUT6), .A3(new_n318), .ZN(new_n319));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n320));
  NOR2_X1   g198(.A1(new_n316), .A2(new_n257), .ZN(new_n321));
  AOI21_X1  g199(.A(new_n321), .B1(new_n276), .B2(new_n125), .ZN(new_n322));
  INV_X1    g200(.A(new_n318), .ZN(new_n323));
  OAI21_X1  g201(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g202(.A1(new_n322), .A2(new_n323), .ZN(new_n325));
  NAND3_X1  g203(.A1(new_n319), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g204(.A1(new_n284), .A2(new_n222), .ZN(new_n327));
  OAI21_X1  g205(.A(new_n327), .B1(new_n222), .B2(new_n162), .ZN(new_n328));
  INV_X1    g206(.A(G224), .ZN(new_n329));
  NOR2_X1   g207(.A1(new_n329), .A2(G953), .ZN(new_n330));
  XNOR2_X1  g208(.A(new_n328), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g209(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g210(.A(new_n328), .B(KEYINPUT7), .C1(new_n329), .C2(G953), .ZN(new_n333));
  INV_X1    g211(.A(KEYINPUT7), .ZN(new_n334));
  OAI221_X1 g212(.A(new_n327), .B1(new_n334), .B2(new_n330), .C1(new_n222), .C2(new_n162), .ZN(new_n335));
  AOI22_X1  g213(.A1(new_n333), .A2(new_n335), .B1(new_n322), .B2(new_n323), .ZN(new_n336));
  XOR2_X1   g214(.A(new_n318), .B(KEYINPUT8), .Z(new_n337));
  AND2_X1   g215(.A1(new_n316), .A2(new_n257), .ZN(new_n338));
  OAI21_X1  g216(.A(new_n337), .B1(new_n338), .B2(new_n321), .ZN(new_n339));
  AOI21_X1  g217(.A(G902), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g218(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n342));
  INV_X1    g220(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g221(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g222(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n345));
  AOI21_X1  g223(.A(new_n307), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g224(.A(G237), .ZN(new_n347));
  NAND3_X1  g225(.A1(new_n347), .A2(new_n227), .A3(G214), .ZN(new_n348));
  NAND2_X1  g226(.A1(new_n348), .A2(new_n135), .ZN(new_n349));
  NAND3_X1  g227(.A1(new_n168), .A2(G143), .A3(G214), .ZN(new_n350));
  NAND2_X1  g228(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g229(.A1(new_n351), .A2(G131), .ZN(new_n352));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g231(.A1(new_n349), .A2(new_n127), .A3(new_n350), .ZN(new_n354));
  NAND3_X1  g232(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g233(.A(new_n218), .ZN(new_n356));
  NAND3_X1  g234(.A1(new_n351), .A2(KEYINPUT17), .A3(G131), .ZN(new_n357));
  NAND4_X1  g235(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(new_n221), .ZN(new_n358));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n359));
  XNOR2_X1  g237(.A(new_n359), .B(new_n251), .ZN(new_n360));
  NAND3_X1  g238(.A1(new_n351), .A2(KEYINPUT18), .A3(G131), .ZN(new_n361));
  XNOR2_X1  g239(.A(new_n212), .B(new_n138), .ZN(new_n362));
  NAND2_X1  g240(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND3_X1  g241(.A1(new_n349), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g242(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g243(.A1(new_n358), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g244(.A1(new_n352), .A2(new_n354), .ZN(new_n367));
  AND2_X1   g245(.A1(new_n212), .A2(KEYINPUT19), .ZN(new_n368));
  NOR2_X1   g246(.A1(new_n212), .A2(KEYINPUT19), .ZN(new_n369));
  OAI21_X1  g247(.A(new_n138), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g248(.A1(new_n367), .A2(new_n221), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g249(.A1(new_n371), .A2(new_n365), .ZN(new_n372));
  OAI21_X1  g250(.A(new_n366), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  INV_X1    g251(.A(G475), .ZN(new_n374));
  NAND3_X1  g252(.A1(new_n373), .A2(new_n374), .A3(new_n197), .ZN(new_n375));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n376));
  NAND2_X1  g254(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g255(.A(new_n366), .ZN(new_n378));
  AOI21_X1  g256(.A(new_n360), .B1(new_n358), .B2(new_n365), .ZN(new_n379));
  OAI21_X1  g257(.A(new_n197), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g258(.A1(new_n380), .A2(G475), .ZN(new_n381));
  NAND4_X1  g259(.A1(new_n373), .A2(KEYINPUT20), .A3(new_n374), .A4(new_n197), .ZN(new_n382));
  NAND3_X1  g260(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n384));
  NAND3_X1  g262(.A1(new_n384), .A2(G952), .A3(new_n227), .ZN(new_n385));
  INV_X1    g263(.A(new_n385), .ZN(new_n386));
  XOR2_X1   g264(.A(KEYINPUT21), .B(G898), .Z(new_n387));
  INV_X1    g265(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g266(.A1(new_n384), .A2(G902), .A3(G953), .ZN(new_n389));
  INV_X1    g267(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g268(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g269(.A(G478), .ZN(new_n392));
  NOR2_X1   g270(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  AOI21_X1  g271(.A(KEYINPUT13), .B1(new_n143), .B2(G143), .ZN(new_n394));
  NOR2_X1   g272(.A1(new_n394), .A2(new_n131), .ZN(new_n395));
  XNOR2_X1  g273(.A(G128), .B(G143), .ZN(new_n396));
  XNOR2_X1  g274(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g275(.A(G116), .B(G122), .ZN(new_n398));
  XNOR2_X1  g276(.A(new_n398), .B(new_n249), .ZN(new_n399));
  NAND2_X1  g277(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g278(.A1(new_n309), .A2(G122), .ZN(new_n401));
  NAND2_X1  g279(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  NAND2_X1  g280(.A1(new_n402), .A2(G107), .ZN(new_n403));
  NAND2_X1  g281(.A1(new_n403), .A2(new_n398), .ZN(new_n404));
  XNOR2_X1  g282(.A(new_n396), .B(new_n131), .ZN(new_n405));
  INV_X1    g283(.A(new_n398), .ZN(new_n406));
  NAND3_X1  g284(.A1(new_n406), .A2(new_n402), .A3(G107), .ZN(new_n407));
  NAND3_X1  g285(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g286(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g287(.A1(new_n244), .A2(new_n234), .A3(G953), .ZN(new_n410));
  INV_X1    g288(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g289(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g290(.A1(new_n400), .A2(new_n408), .A3(new_n410), .ZN(new_n413));
  NAND2_X1  g291(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g292(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g293(.A(new_n393), .B1(new_n415), .B2(G902), .ZN(new_n416));
  OAI211_X1 g294(.A(new_n414), .B(new_n197), .C1(KEYINPUT15), .C2(new_n392), .ZN(new_n417));
  NAND2_X1  g295(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR3_X1   g296(.A1(new_n383), .A2(new_n391), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g297(.A1(new_n346), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g298(.A1(new_n305), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g299(.A(new_n421), .B(new_n247), .ZN(G3));
  NAND2_X1  g300(.A1(new_n414), .A2(KEYINPUT33), .ZN(new_n423));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n424));
  NAND3_X1  g302(.A1(new_n412), .A2(new_n424), .A3(new_n413), .ZN(new_n425));
  NAND3_X1  g303(.A1(new_n423), .A2(G478), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g304(.A1(new_n414), .A2(new_n392), .A3(new_n197), .ZN(new_n427));
  NAND2_X1  g305(.A1(G478), .A2(G902), .ZN(new_n428));
  NAND3_X1  g306(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g307(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g308(.A1(new_n430), .A2(new_n383), .ZN(new_n431));
  INV_X1    g309(.A(new_n431), .ZN(new_n432));
  INV_X1    g310(.A(new_n391), .ZN(new_n433));
  NAND3_X1  g311(.A1(new_n432), .A2(new_n346), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g312(.A1(new_n188), .A2(new_n197), .ZN(new_n435));
  AOI22_X1  g313(.A1(new_n435), .A2(G472), .B1(new_n189), .B2(new_n188), .ZN(new_n436));
  NAND3_X1  g314(.A1(new_n304), .A2(new_n436), .A3(new_n243), .ZN(new_n437));
  NOR2_X1   g315(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g316(.A(KEYINPUT34), .B(G104), .ZN(new_n439));
  XNOR2_X1  g317(.A(new_n438), .B(new_n439), .ZN(G6));
  AOI21_X1  g318(.A(new_n383), .B1(new_n417), .B2(new_n416), .ZN(new_n441));
  NAND3_X1  g319(.A1(new_n346), .A2(new_n441), .A3(new_n433), .ZN(new_n442));
  NOR2_X1   g320(.A1(new_n442), .A2(new_n437), .ZN(new_n443));
  XNOR2_X1  g321(.A(KEYINPUT35), .B(G107), .ZN(new_n444));
  XNOR2_X1  g322(.A(new_n443), .B(new_n444), .ZN(G9));
  NAND3_X1  g323(.A1(new_n346), .A2(new_n304), .A3(new_n419), .ZN(new_n446));
  NAND2_X1  g324(.A1(new_n219), .A2(new_n225), .ZN(new_n447));
  NOR2_X1   g325(.A1(new_n229), .A2(KEYINPUT36), .ZN(new_n448));
  XNOR2_X1  g326(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g327(.A1(new_n449), .A2(new_n240), .ZN(new_n450));
  AND2_X1   g328(.A1(new_n238), .A2(new_n450), .ZN(new_n451));
  INV_X1    g329(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g330(.A1(new_n436), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g331(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g332(.A(KEYINPUT37), .B(G110), .ZN(new_n455));
  XNOR2_X1  g333(.A(new_n454), .B(new_n455), .ZN(G12));
  NAND4_X1  g334(.A1(new_n202), .A2(new_n304), .A3(new_n346), .A4(new_n452), .ZN(new_n457));
  INV_X1    g335(.A(G900), .ZN(new_n458));
  AOI21_X1  g336(.A(new_n386), .B1(new_n390), .B2(new_n458), .ZN(new_n459));
  INV_X1    g337(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g338(.A1(new_n441), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g339(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g340(.A(new_n462), .B(new_n143), .ZN(G30));
  XOR2_X1   g341(.A(new_n459), .B(KEYINPUT39), .Z(new_n464));
  NAND2_X1  g342(.A1(new_n304), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g343(.A(new_n465), .B(KEYINPUT40), .Z(new_n466));
  AND3_X1   g344(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n467));
  AOI21_X1  g345(.A(new_n342), .B1(new_n332), .B2(new_n340), .ZN(new_n468));
  NOR2_X1   g346(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g347(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n470));
  NAND2_X1  g348(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n471));
  NAND2_X1  g349(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g350(.A1(new_n472), .A2(new_n452), .ZN(new_n473));
  AND2_X1   g351(.A1(new_n184), .A2(new_n167), .ZN(new_n474));
  NOR2_X1   g352(.A1(new_n474), .A2(new_n180), .ZN(new_n475));
  NAND3_X1  g353(.A1(new_n177), .A2(new_n180), .A3(new_n167), .ZN(new_n476));
  NAND2_X1  g354(.A1(new_n476), .A2(new_n197), .ZN(new_n477));
  OAI21_X1  g355(.A(G472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g356(.A1(new_n192), .A2(new_n201), .A3(new_n478), .ZN(new_n479));
  INV_X1    g357(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g358(.A1(new_n383), .A2(new_n418), .ZN(new_n481));
  NOR2_X1   g359(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g360(.A1(new_n466), .A2(new_n473), .A3(new_n306), .A4(new_n482), .ZN(new_n483));
  XNOR2_X1  g361(.A(new_n483), .B(G143), .ZN(G45));
  NOR2_X1   g362(.A1(new_n431), .A2(new_n459), .ZN(new_n485));
  INV_X1    g363(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g364(.A1(new_n457), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g365(.A(new_n487), .B(new_n138), .ZN(G48));
  OAI21_X1  g366(.A(new_n197), .B1(new_n301), .B2(new_n302), .ZN(new_n489));
  NAND2_X1  g367(.A1(new_n489), .A2(G469), .ZN(new_n490));
  AND3_X1   g368(.A1(new_n490), .A2(new_n245), .A3(new_n303), .ZN(new_n491));
  NAND3_X1  g369(.A1(new_n202), .A2(new_n243), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g370(.A1(new_n492), .A2(new_n434), .ZN(new_n493));
  XOR2_X1   g371(.A(KEYINPUT41), .B(G113), .Z(new_n494));
  XNOR2_X1  g372(.A(new_n493), .B(new_n494), .ZN(G15));
  NOR2_X1   g373(.A1(new_n492), .A2(new_n442), .ZN(new_n496));
  XNOR2_X1  g374(.A(new_n496), .B(new_n309), .ZN(G18));
  NOR2_X1   g375(.A1(new_n383), .A2(new_n418), .ZN(new_n498));
  NAND3_X1  g376(.A1(new_n202), .A2(new_n498), .A3(new_n452), .ZN(new_n499));
  NAND3_X1  g377(.A1(new_n491), .A2(new_n346), .A3(new_n433), .ZN(new_n500));
  NOR2_X1   g378(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g379(.A(new_n501), .B(new_n204), .ZN(G21));
  NAND4_X1  g380(.A1(new_n436), .A2(new_n243), .A3(new_n383), .A4(new_n418), .ZN(new_n503));
  NOR2_X1   g381(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g382(.A(new_n504), .B(G122), .Z(G24));
  INV_X1    g383(.A(new_n190), .ZN(new_n506));
  INV_X1    g384(.A(G472), .ZN(new_n507));
  AOI21_X1  g385(.A(new_n507), .B1(new_n188), .B2(new_n197), .ZN(new_n508));
  NOR3_X1   g386(.A1(new_n506), .A2(new_n508), .A3(new_n451), .ZN(new_n509));
  NAND4_X1  g387(.A1(new_n509), .A2(new_n485), .A3(new_n346), .A4(new_n491), .ZN(new_n510));
  XNOR2_X1  g388(.A(new_n510), .B(G125), .ZN(G27));
  NOR3_X1   g389(.A1(new_n467), .A2(new_n468), .A3(new_n307), .ZN(new_n512));
  AND4_X1   g390(.A1(new_n202), .A2(new_n243), .A3(new_n304), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g391(.A1(new_n513), .A2(KEYINPUT42), .A3(new_n485), .ZN(new_n514));
  INV_X1    g392(.A(KEYINPUT42), .ZN(new_n515));
  NAND4_X1  g393(.A1(new_n202), .A2(new_n243), .A3(new_n304), .A4(new_n512), .ZN(new_n516));
  OAI21_X1  g394(.A(new_n515), .B1(new_n516), .B2(new_n486), .ZN(new_n517));
  NAND2_X1  g395(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g396(.A(new_n518), .B(G131), .ZN(G33));
  NOR2_X1   g397(.A1(new_n516), .A2(new_n461), .ZN(new_n520));
  XNOR2_X1  g398(.A(new_n520), .B(new_n131), .ZN(G36));
  NAND2_X1  g399(.A1(new_n291), .A2(KEYINPUT45), .ZN(new_n522));
  INV_X1    g400(.A(KEYINPUT45), .ZN(new_n523));
  NAND3_X1  g401(.A1(new_n271), .A2(new_n278), .A3(new_n282), .ZN(new_n524));
  INV_X1    g402(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g403(.A(new_n282), .B1(new_n300), .B2(new_n278), .ZN(new_n526));
  OAI21_X1  g404(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g405(.A1(new_n522), .A2(G469), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g406(.A1(G469), .A2(G902), .ZN(new_n529));
  NAND3_X1  g407(.A1(new_n528), .A2(KEYINPUT46), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g408(.A1(new_n530), .A2(new_n303), .ZN(new_n531));
  AOI21_X1  g409(.A(KEYINPUT46), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  OAI211_X1 g410(.A(new_n245), .B(new_n464), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n534));
  INV_X1    g412(.A(new_n436), .ZN(new_n535));
  OR3_X1    g413(.A1(new_n383), .A2(new_n429), .A3(KEYINPUT43), .ZN(new_n536));
  OAI21_X1  g414(.A(KEYINPUT43), .B1(new_n383), .B2(new_n429), .ZN(new_n537));
  NAND4_X1  g415(.A1(new_n535), .A2(new_n536), .A3(new_n452), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g416(.A(new_n533), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g417(.A1(new_n538), .A2(new_n534), .ZN(new_n540));
  INV_X1    g418(.A(new_n512), .ZN(new_n541));
  NOR2_X1   g419(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g420(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g421(.A(new_n543), .B(G137), .ZN(G39));
  OAI21_X1  g422(.A(new_n245), .B1(new_n531), .B2(new_n532), .ZN(new_n545));
  INV_X1    g423(.A(KEYINPUT47), .ZN(new_n546));
  NAND2_X1  g424(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g425(.A(KEYINPUT47), .B(new_n245), .C1(new_n531), .C2(new_n532), .ZN(new_n548));
  NAND2_X1  g426(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g427(.A1(new_n541), .A2(new_n202), .A3(new_n243), .ZN(new_n550));
  NAND3_X1  g428(.A1(new_n549), .A2(new_n485), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g429(.A(new_n551), .B(G140), .ZN(G42));
  AND3_X1   g430(.A1(new_n536), .A2(new_n386), .A3(new_n537), .ZN(new_n553));
  NOR2_X1   g431(.A1(new_n535), .A2(new_n242), .ZN(new_n554));
  AND2_X1   g432(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g433(.A1(new_n490), .A2(new_n303), .ZN(new_n556));
  AND2_X1   g434(.A1(new_n556), .A2(new_n246), .ZN(new_n557));
  OAI211_X1 g435(.A(new_n512), .B(new_n555), .C1(new_n549), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g436(.A(new_n306), .B1(new_n470), .B2(new_n471), .ZN(new_n559));
  NAND4_X1  g437(.A1(new_n555), .A2(KEYINPUT50), .A3(new_n491), .A4(new_n559), .ZN(new_n560));
  INV_X1    g438(.A(KEYINPUT50), .ZN(new_n561));
  INV_X1    g439(.A(new_n559), .ZN(new_n562));
  NAND3_X1  g440(.A1(new_n553), .A2(new_n554), .A3(new_n491), .ZN(new_n563));
  OAI21_X1  g441(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g442(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g443(.A1(new_n491), .A2(new_n512), .ZN(new_n566));
  NAND2_X1  g444(.A1(new_n480), .A2(new_n386), .ZN(new_n567));
  NOR4_X1   g445(.A1(new_n567), .A2(new_n242), .A3(new_n383), .A4(new_n430), .ZN(new_n568));
  AND2_X1   g446(.A1(new_n553), .A2(new_n509), .ZN(new_n569));
  OAI21_X1  g447(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g448(.A1(new_n558), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g449(.A(new_n571), .B(KEYINPUT51), .ZN(new_n572));
  INV_X1    g450(.A(G952), .ZN(new_n573));
  NOR3_X1   g451(.A1(new_n567), .A2(new_n242), .A3(new_n431), .ZN(new_n574));
  AOI211_X1 g452(.A(new_n573), .B(G953), .C1(new_n574), .C2(new_n566), .ZN(new_n575));
  AND2_X1   g453(.A1(new_n202), .A2(new_n243), .ZN(new_n576));
  NAND3_X1  g454(.A1(new_n553), .A2(new_n576), .A3(new_n566), .ZN(new_n577));
  XNOR2_X1  g455(.A(new_n577), .B(KEYINPUT48), .ZN(new_n578));
  NAND3_X1  g456(.A1(new_n555), .A2(new_n346), .A3(new_n491), .ZN(new_n579));
  AND3_X1   g457(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND4_X1   g458(.A1(new_n202), .A2(new_n304), .A3(new_n346), .A4(new_n452), .ZN(new_n581));
  INV_X1    g459(.A(new_n461), .ZN(new_n582));
  OAI21_X1  g460(.A(new_n581), .B1(new_n582), .B2(new_n485), .ZN(new_n583));
  INV_X1    g461(.A(KEYINPUT52), .ZN(new_n584));
  OAI21_X1  g462(.A(new_n306), .B1(new_n467), .B2(new_n468), .ZN(new_n585));
  NOR2_X1   g463(.A1(new_n585), .A2(new_n481), .ZN(new_n586));
  NAND2_X1  g464(.A1(new_n289), .A2(new_n290), .ZN(new_n587));
  NAND3_X1  g465(.A1(new_n587), .A2(G469), .A3(new_n524), .ZN(new_n588));
  NAND3_X1  g466(.A1(new_n303), .A2(new_n529), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g467(.A1(new_n589), .A2(new_n245), .A3(new_n460), .ZN(new_n590));
  NAND4_X1  g468(.A1(new_n586), .A2(new_n451), .A3(new_n479), .A4(new_n590), .ZN(new_n591));
  NAND4_X1  g469(.A1(new_n583), .A2(new_n584), .A3(new_n510), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g470(.A(new_n457), .B1(new_n461), .B2(new_n486), .ZN(new_n593));
  NAND2_X1  g471(.A1(new_n591), .A2(new_n510), .ZN(new_n594));
  OAI21_X1  g472(.A(KEYINPUT52), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g473(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g474(.A(new_n520), .ZN(new_n597));
  NAND3_X1  g475(.A1(new_n432), .A2(new_n436), .A3(new_n452), .ZN(new_n598));
  NAND2_X1  g476(.A1(new_n499), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g477(.A1(new_n599), .A2(new_n512), .A3(new_n590), .ZN(new_n600));
  AOI21_X1  g478(.A(KEYINPUT42), .B1(new_n513), .B2(new_n485), .ZN(new_n601));
  NOR3_X1   g479(.A1(new_n516), .A2(new_n515), .A3(new_n486), .ZN(new_n602));
  OAI211_X1 g480(.A(new_n597), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g481(.A(new_n603), .ZN(new_n604));
  OAI22_X1  g482(.A1(new_n492), .A2(new_n434), .B1(new_n500), .B2(new_n503), .ZN(new_n605));
  NOR2_X1   g483(.A1(new_n605), .A2(new_n496), .ZN(new_n606));
  OAI22_X1  g484(.A1(new_n305), .A2(new_n420), .B1(new_n446), .B2(new_n453), .ZN(new_n607));
  AOI21_X1  g485(.A(new_n437), .B1(new_n434), .B2(new_n442), .ZN(new_n608));
  NOR2_X1   g486(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g487(.A(new_n501), .ZN(new_n610));
  AND3_X1   g488(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g489(.A1(new_n596), .A2(KEYINPUT53), .A3(new_n604), .A4(new_n611), .ZN(new_n612));
  INV_X1    g490(.A(KEYINPUT53), .ZN(new_n613));
  NOR3_X1   g491(.A1(new_n607), .A2(new_n608), .A3(new_n501), .ZN(new_n614));
  INV_X1    g492(.A(new_n590), .ZN(new_n615));
  AOI21_X1  g493(.A(new_n615), .B1(new_n499), .B2(new_n598), .ZN(new_n616));
  AOI21_X1  g494(.A(new_n520), .B1(new_n512), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g495(.A1(new_n614), .A2(new_n617), .A3(new_n518), .A4(new_n606), .ZN(new_n618));
  NAND2_X1  g496(.A1(new_n592), .A2(new_n595), .ZN(new_n619));
  OAI21_X1  g497(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g498(.A(KEYINPUT54), .B1(new_n612), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g499(.A1(new_n612), .A2(KEYINPUT54), .A3(new_n620), .ZN(new_n622));
  OAI211_X1 g500(.A(new_n572), .B(new_n580), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g501(.A1(new_n573), .A2(new_n227), .ZN(new_n624));
  NAND2_X1  g502(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g503(.A(new_n556), .B(KEYINPUT49), .Z(new_n626));
  NOR2_X1   g504(.A1(new_n626), .A2(new_n479), .ZN(new_n627));
  NOR2_X1   g505(.A1(new_n383), .A2(new_n429), .ZN(new_n628));
  NOR3_X1   g506(.A1(new_n242), .A2(new_n246), .A3(new_n307), .ZN(new_n629));
  NAND4_X1  g507(.A1(new_n627), .A2(new_n472), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g508(.A1(new_n625), .A2(new_n630), .ZN(G75));
  NAND2_X1  g509(.A1(new_n612), .A2(new_n620), .ZN(new_n632));
  NAND3_X1  g510(.A1(new_n632), .A2(G902), .A3(new_n343), .ZN(new_n633));
  INV_X1    g511(.A(KEYINPUT56), .ZN(new_n634));
  XOR2_X1   g512(.A(new_n326), .B(new_n331), .Z(new_n635));
  XNOR2_X1  g513(.A(new_n635), .B(KEYINPUT55), .ZN(new_n636));
  AND3_X1   g514(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g515(.A(new_n636), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  NOR2_X1   g516(.A1(new_n227), .A2(G952), .ZN(new_n639));
  NOR3_X1   g517(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(G51));
  INV_X1    g518(.A(KEYINPUT54), .ZN(new_n641));
  NAND3_X1  g519(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n642));
  NOR2_X1   g520(.A1(new_n642), .A2(new_n603), .ZN(new_n643));
  AOI21_X1  g521(.A(KEYINPUT53), .B1(new_n643), .B2(new_n596), .ZN(new_n644));
  NOR3_X1   g522(.A1(new_n618), .A2(new_n619), .A3(new_n613), .ZN(new_n645));
  OAI21_X1  g523(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g524(.A1(new_n612), .A2(KEYINPUT54), .A3(new_n620), .ZN(new_n647));
  XOR2_X1   g525(.A(new_n529), .B(KEYINPUT57), .Z(new_n648));
  NAND3_X1  g526(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g527(.A1(new_n301), .A2(new_n302), .ZN(new_n650));
  NAND2_X1  g528(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g529(.A(new_n528), .ZN(new_n652));
  NAND3_X1  g530(.A1(new_n632), .A2(G902), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g531(.A(new_n639), .B1(new_n651), .B2(new_n653), .ZN(G54));
  AND2_X1   g532(.A1(new_n632), .A2(KEYINPUT58), .ZN(new_n655));
  NOR2_X1   g533(.A1(new_n374), .A2(new_n197), .ZN(new_n656));
  AOI21_X1  g534(.A(new_n373), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g535(.A1(new_n632), .A2(KEYINPUT58), .A3(new_n373), .A4(new_n656), .ZN(new_n658));
  INV_X1    g536(.A(new_n639), .ZN(new_n659));
  NAND2_X1  g537(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g538(.A1(new_n657), .A2(new_n660), .ZN(G60));
  XNOR2_X1  g539(.A(new_n428), .B(KEYINPUT59), .ZN(new_n662));
  NAND3_X1  g540(.A1(new_n646), .A2(new_n647), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g541(.A1(new_n423), .A2(new_n425), .ZN(new_n664));
  INV_X1    g542(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g543(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g544(.A1(new_n646), .A2(new_n664), .A3(new_n647), .A4(new_n662), .ZN(new_n667));
  AND3_X1   g545(.A1(new_n666), .A2(new_n659), .A3(new_n667), .ZN(G63));
  INV_X1    g546(.A(KEYINPUT61), .ZN(new_n669));
  NAND2_X1  g547(.A1(G217), .A2(G902), .ZN(new_n670));
  XOR2_X1   g548(.A(new_n670), .B(KEYINPUT60), .Z(new_n671));
  NAND3_X1  g549(.A1(new_n632), .A2(new_n449), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g550(.A1(new_n672), .A2(new_n659), .ZN(new_n673));
  AOI21_X1  g551(.A(new_n239), .B1(new_n632), .B2(new_n671), .ZN(new_n674));
  OAI21_X1  g552(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g553(.A(new_n674), .ZN(new_n676));
  NAND4_X1  g554(.A1(new_n676), .A2(KEYINPUT61), .A3(new_n659), .A4(new_n672), .ZN(new_n677));
  NAND2_X1  g555(.A1(new_n675), .A2(new_n677), .ZN(G66));
  OAI21_X1  g556(.A(G953), .B1(new_n388), .B2(new_n329), .ZN(new_n679));
  OAI21_X1  g557(.A(new_n679), .B1(new_n611), .B2(G953), .ZN(new_n680));
  INV_X1    g558(.A(new_n326), .ZN(new_n681));
  OAI21_X1  g559(.A(new_n681), .B1(G898), .B2(new_n227), .ZN(new_n682));
  XNOR2_X1  g560(.A(new_n680), .B(new_n682), .ZN(G69));
  NAND2_X1  g561(.A1(new_n161), .A2(new_n165), .ZN(new_n684));
  NOR2_X1   g562(.A1(new_n368), .A2(new_n369), .ZN(new_n685));
  XOR2_X1   g563(.A(new_n684), .B(new_n685), .Z(new_n686));
  OAI21_X1  g564(.A(new_n686), .B1(G900), .B2(new_n227), .ZN(new_n687));
  OAI21_X1  g565(.A(G953), .B1(new_n280), .B2(new_n458), .ZN(new_n688));
  NOR2_X1   g566(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g567(.A1(new_n483), .A2(new_n510), .A3(new_n583), .ZN(new_n690));
  NAND2_X1  g568(.A1(new_n690), .A2(KEYINPUT62), .ZN(new_n691));
  AND2_X1   g569(.A1(new_n551), .A2(new_n543), .ZN(new_n692));
  INV_X1    g570(.A(KEYINPUT62), .ZN(new_n693));
  NAND4_X1  g571(.A1(new_n483), .A2(new_n693), .A3(new_n510), .A4(new_n583), .ZN(new_n694));
  NOR2_X1   g572(.A1(new_n465), .A2(new_n541), .ZN(new_n695));
  OAI211_X1 g573(.A(new_n695), .B(new_n576), .C1(new_n432), .C2(new_n441), .ZN(new_n696));
  NAND4_X1  g574(.A1(new_n691), .A2(new_n692), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g575(.A1(new_n697), .A2(new_n227), .ZN(new_n698));
  NAND2_X1  g576(.A1(new_n698), .A2(new_n687), .ZN(new_n699));
  AND3_X1   g577(.A1(new_n543), .A2(new_n510), .A3(new_n597), .ZN(new_n700));
  NAND2_X1  g578(.A1(new_n576), .A2(new_n586), .ZN(new_n701));
  NOR2_X1   g579(.A1(new_n533), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g580(.A1(new_n702), .A2(new_n593), .ZN(new_n703));
  NAND4_X1  g581(.A1(new_n700), .A2(new_n518), .A3(new_n551), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g582(.A1(new_n704), .A2(new_n227), .A3(new_n686), .ZN(new_n705));
  NAND2_X1  g583(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g584(.A(new_n689), .B1(new_n706), .B2(new_n688), .ZN(G72));
  NAND2_X1  g585(.A1(G472), .A2(G902), .ZN(new_n708));
  XOR2_X1   g586(.A(new_n708), .B(KEYINPUT63), .Z(new_n709));
  OAI21_X1  g587(.A(new_n709), .B1(new_n704), .B2(new_n642), .ZN(new_n710));
  NAND2_X1  g588(.A1(new_n474), .A2(new_n180), .ZN(new_n711));
  INV_X1    g589(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g590(.A(new_n639), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g591(.A(new_n709), .B1(new_n697), .B2(new_n642), .ZN(new_n714));
  NAND2_X1  g592(.A1(new_n714), .A2(new_n475), .ZN(new_n715));
  INV_X1    g593(.A(new_n475), .ZN(new_n716));
  NAND4_X1  g594(.A1(new_n632), .A2(new_n716), .A3(new_n709), .A4(new_n711), .ZN(new_n717));
  AND3_X1   g595(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(G57));
endmodule


