//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(KEYINPUT66), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(KEYINPUT66), .B2(new_n457), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n460), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n461), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(new_n465), .B(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n476), .A2(G136), .B1(G124), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND3_X1  g058(.A1(new_n471), .A2(G138), .A3(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n465), .A2(G138), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n491), .B1(new_n490), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n489), .B(new_n498), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n504), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n518), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n505), .A2(new_n514), .A3(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND3_X1  g103(.A1(new_n502), .A2(new_n504), .A3(G64), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n532), .A2(G651), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT73), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n516), .A2(G90), .B1(G52), .B2(new_n518), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n532), .A2(new_n538), .A3(G651), .A4(new_n534), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  XOR2_X1   g116(.A(KEYINPUT75), .B(G81), .Z(new_n542));
  AOI22_X1  g117(.A1(new_n516), .A2(new_n542), .B1(new_n518), .B2(G43), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  INV_X1    g119(.A(G68), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n509), .A2(new_n544), .B1(new_n545), .B2(new_n501), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI221_X1 g123(.A(KEYINPUT74), .B1(new_n545), .B2(new_n501), .C1(new_n509), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n509), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n516), .A2(G91), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G299));
  NAND2_X1  g140(.A1(new_n516), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n518), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G651), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n515), .A2(new_n573), .B1(new_n517), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n516), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n578));
  NAND2_X1  g153(.A1(G72), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G60), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n509), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G290));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n509), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(G54), .A2(new_n518), .B1(new_n588), .B2(G651), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT10), .B1(new_n515), .B2(new_n584), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G171), .B2(new_n592), .ZN(G321));
  XOR2_X1   g169(.A(G321), .B(KEYINPUT76), .Z(G284));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(new_n591), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n551), .A2(new_n592), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n591), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n592), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n476), .A2(G135), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n478), .A2(G123), .ZN(new_n609));
  OR2_X1    g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2096), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n471), .A2(new_n467), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XOR2_X1   g191(.A(KEYINPUT13), .B(G2100), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2430), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XOR2_X1   g200(.A(G2443), .B(G2446), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G14), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XOR2_X1   g210(.A(G2072), .B(G2078), .Z(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT80), .Z(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n637), .B(KEYINPUT17), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n641), .B2(new_n638), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(new_n643));
  INV_X1    g218(.A(new_n637), .ZN(new_n644));
  INV_X1    g219(.A(new_n638), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(new_n635), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT18), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n638), .A3(new_n635), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n654), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT84), .B(G1981), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n670), .B(new_n673), .Z(G229));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(G28), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(G28), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n676), .A2(new_n677), .A3(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(G171), .A2(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G5), .B2(G16), .ZN(new_n680));
  INV_X1    g255(.A(G1961), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(KEYINPUT91), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT31), .B(G11), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(G16), .A2(G21), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G168), .B2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G1966), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n612), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n687), .A2(KEYINPUT92), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n685), .A2(new_n691), .A3(new_n693), .A4(new_n686), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(KEYINPUT23), .A3(G20), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT23), .ZN(new_n700));
  INV_X1    g275(.A(G20), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G16), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n702), .C1(new_n597), .C2(new_n698), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1956), .ZN(new_n704));
  INV_X1    g279(.A(G1348), .ZN(new_n705));
  NOR2_X1   g280(.A1(G4), .A2(G16), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n600), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n704), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n692), .A2(G26), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n476), .A2(G140), .B1(G128), .B2(new_n478), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT88), .B(G2067), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT24), .A2(G34), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(new_n692), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G160), .B2(new_n692), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G32), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n467), .A2(G105), .ZN(new_n731));
  INV_X1    g306(.A(G129), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n477), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n476), .B2(G141), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n709), .A2(new_n721), .A3(new_n727), .A4(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n692), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n482), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n692), .A2(G33), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT90), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n467), .A2(G103), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n476), .A2(G139), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n748), .B(new_n749), .C1(new_n470), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n744), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G2072), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n680), .A2(new_n681), .B1(G1348), .B2(new_n707), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n743), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(new_n720), .B2(new_n718), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n738), .A2(new_n757), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n694), .A2(new_n697), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n741), .A2(new_n742), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n698), .A2(G22), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G166), .B2(new_n698), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1971), .ZN(new_n770));
  NOR2_X1   g345(.A1(G6), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n576), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT32), .B(G1981), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(G1971), .ZN(new_n775));
  OR2_X1    g350(.A1(G16), .A2(G23), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G288), .B2(new_n698), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT33), .B(G1976), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n770), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT85), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT85), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT86), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(KEYINPUT86), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n476), .A2(G131), .B1(G119), .B2(new_n478), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n470), .A2(G107), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n698), .A2(G24), .ZN(new_n798));
  INV_X1    g373(.A(G290), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n698), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(new_n667), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n796), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n767), .B1(new_n789), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g379(.A(KEYINPUT36), .B(new_n802), .C1(new_n787), .C2(new_n788), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n765), .B(new_n766), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n698), .A2(G19), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n552), .B2(new_n698), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1341), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT93), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n694), .A2(new_n697), .A3(new_n764), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n789), .A2(new_n803), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n789), .A2(new_n767), .A3(new_n803), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n816));
  INV_X1    g391(.A(new_n809), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n766), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n810), .A2(new_n818), .ZN(G311));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n766), .A3(new_n817), .ZN(G150));
  AOI22_X1  g395(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n571), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n518), .A2(G55), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n505), .A2(new_n514), .A3(G93), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n823), .A2(KEYINPUT94), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT94), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n551), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n601), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n834), .B2(G860), .ZN(G145));
  INV_X1    g410(.A(G37), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n482), .B(KEYINPUT95), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G160), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n612), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n717), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n490), .A2(new_n493), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n489), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n734), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n842), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT97), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT97), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n849), .B(new_n850), .C1(G118), .C2(new_n470), .ZN(new_n851));
  INV_X1    g426(.A(G130), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n477), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n476), .B2(G142), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n616), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n793), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n847), .A2(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n840), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n857), .A2(new_n860), .A3(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n839), .B1(new_n857), .B2(new_n860), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n836), .B(new_n859), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(new_n827), .A2(new_n592), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n827), .B(new_n552), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n604), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(G299), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT99), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n591), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n600), .A2(new_n597), .A3(KEYINPUT99), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT41), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(new_n872), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n866), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n866), .B2(new_n881), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G288), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT101), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(new_n576), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n886), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n887), .A2(KEYINPUT42), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(new_n890), .C1(new_n885), .C2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n892), .B1(new_n896), .B2(KEYINPUT42), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n883), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n865), .B1(new_n898), .B2(new_n592), .ZN(G295));
  OAI21_X1  g474(.A(new_n865), .B1(new_n898), .B2(new_n592), .ZN(G331));
  NAND2_X1  g475(.A1(G301), .A2(G168), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND3_X1  g478(.A1(G301), .A2(new_n903), .A3(G168), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n536), .A2(G286), .A3(new_n537), .A4(new_n539), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT104), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n905), .A2(new_n830), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n830), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n876), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  AND3_X1   g486(.A1(G301), .A2(new_n903), .A3(G168), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n903), .B1(G301), .B2(G168), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n906), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n867), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n905), .A2(new_n907), .A3(new_n830), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n876), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n905), .A2(new_n907), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n867), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n908), .A2(new_n909), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n926), .B(new_n880), .C1(new_n927), .C2(KEYINPUT106), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n896), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT107), .B1(new_n929), .B2(G37), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n923), .B2(new_n919), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n911), .A2(new_n921), .B1(new_n931), .B2(new_n880), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n896), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n836), .C1(new_n932), .C2(new_n896), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n919), .A2(new_n879), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n926), .B1(new_n927), .B2(KEYINPUT106), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n876), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n896), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT108), .B1(new_n941), .B2(new_n896), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(KEYINPUT43), .A3(new_n933), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n944), .A2(new_n937), .A3(new_n933), .A4(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(G397));
  AND2_X1   g529(.A1(G160), .A2(G40), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n845), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G1996), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT110), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n959), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n717), .B(G2067), .Z(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n734), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n962), .A2(new_n734), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n793), .B(new_n795), .Z(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(G1986), .A3(G290), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n667), .A3(new_n799), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT109), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(G301), .B(KEYINPUT54), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n843), .B1(new_n488), .B2(new_n487), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n978), .B2(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n845), .A2(KEYINPUT111), .A3(new_n957), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n497), .A2(new_n957), .A3(new_n499), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT122), .B(G1961), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n955), .B1(new_n958), .B2(new_n956), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n984), .B2(new_n956), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n760), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n991), .A2(KEYINPUT123), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT123), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n957), .A4(new_n499), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n979), .A2(new_n980), .A3(new_n956), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n955), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n998), .A2(new_n992), .A3(G2078), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n983), .A2(new_n726), .A3(new_n985), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n690), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1009), .A2(KEYINPUT121), .B1(new_n1008), .B2(G168), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G168), .A2(new_n1008), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(KEYINPUT120), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(KEYINPUT120), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1007), .A2(new_n1010), .B1(new_n1015), .B2(new_n1001), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n975), .A2(new_n1000), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n984), .A2(new_n956), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n989), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n986), .B2(G2090), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(G8), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n1008), .ZN(new_n1028));
  INV_X1    g603(.A(G288), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G1976), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n576), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n572), .B2(new_n575), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1033), .B(KEYINPUT49), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(new_n1027), .A3(new_n1008), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT49), .B1(new_n1039), .B2(new_n1033), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1028), .A2(new_n1030), .A3(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1032), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1026), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT124), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n474), .B1(new_n469), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(G40), .C1(new_n1047), .C2(new_n469), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT125), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n958), .A2(new_n956), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n958), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1051), .B(new_n1054), .C1(KEYINPUT45), .C2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n992), .A2(G2078), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n975), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n988), .C1(new_n993), .C2(new_n994), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT50), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n955), .C1(new_n984), .C2(KEYINPUT50), .ZN(new_n1061));
  OAI22_X1  g636(.A1(G1971), .A2(new_n990), .B1(new_n1061), .B2(G2090), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1025), .B1(new_n1062), .B2(G8), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1046), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1018), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n990), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(G299), .B(KEYINPUT57), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n990), .A2(new_n965), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1027), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n552), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  OAI221_X1 g661(.A(new_n552), .B1(KEYINPUT116), .B2(new_n1086), .C1(new_n1078), .C2(new_n1082), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1075), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n1089));
  OR2_X1    g664(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1090), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1073), .A2(KEYINPUT118), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n986), .A2(new_n705), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1079), .A2(G2067), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n983), .B2(new_n985), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT114), .B1(new_n1104), .B2(new_n1100), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n600), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1102), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1104), .A2(new_n1100), .A3(KEYINPUT114), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT119), .A3(new_n591), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1108), .A2(new_n1112), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1088), .B(new_n1097), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1114), .A2(new_n1092), .A3(new_n591), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1091), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1066), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1000), .A2(new_n1064), .A3(new_n1046), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1016), .A2(KEYINPUT62), .A3(new_n1017), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT62), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1120), .B(G171), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1009), .A2(new_n1124), .A3(G168), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1026), .B1(new_n1125), .B2(new_n1063), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1126), .A2(new_n1045), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1021), .B(new_n1024), .C1(new_n986), .C2(G2090), .ZN(new_n1128));
  AOI22_X1  g703(.A1(KEYINPUT52), .A2(new_n1031), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1044), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1009), .A2(G168), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT63), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1041), .A2(new_n1042), .A3(new_n1029), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1035), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1028), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT113), .B1(new_n1127), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1126), .A2(new_n1045), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(new_n1135), .A4(new_n1132), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1123), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n974), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n717), .A2(G2067), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n793), .A2(new_n795), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n967), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n959), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT126), .Z(new_n1148));
  XOR2_X1   g723(.A(new_n971), .B(KEYINPUT48), .Z(new_n1149));
  NOR2_X1   g724(.A1(new_n969), .A2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n964), .A2(new_n734), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1151), .A2(new_n1152), .B1(new_n959), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1155));
  XNOR2_X1  g730(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1148), .A2(new_n1150), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g733(.A1(G319), .A2(new_n863), .A3(new_n633), .A4(new_n651), .ZN(new_n1160));
  INV_X1    g734(.A(G229), .ZN(new_n1161));
  AND3_X1   g735(.A1(new_n1160), .A2(new_n951), .A3(new_n1161), .ZN(G308));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n951), .A3(new_n1161), .ZN(G225));
endmodule


