//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  OAI211_X1 g002(.A(new_n187), .B(G146), .C1(new_n188), .C2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT66), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n197), .A3(new_n191), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT80), .A2(G104), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT80), .A2(G104), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(KEYINPUT81), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n207), .A3(new_n201), .A4(new_n202), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G101), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(new_n202), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n204), .A2(KEYINPUT3), .A3(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n215), .A3(KEYINPUT84), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n199), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n216), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n192), .A2(KEYINPUT82), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n192), .A2(KEYINPUT82), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n196), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G134), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT11), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n227), .A3(G134), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(G137), .ZN(new_n237));
  AND4_X1   g051(.A1(KEYINPUT64), .A2(new_n236), .A3(new_n234), .A4(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT64), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT12), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n241), .A2(KEYINPUT12), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n226), .A2(new_n240), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n220), .A2(new_n225), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n233), .A2(new_n234), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n231), .B1(G134), .B2(new_n227), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n229), .A2(KEYINPUT11), .A3(G137), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n234), .B(new_n237), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n233), .A2(KEYINPUT64), .A3(new_n234), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n241), .B(KEYINPUT12), .C1(new_n245), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n221), .A2(new_n224), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n218), .A2(KEYINPUT10), .A3(new_n199), .A4(new_n219), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n194), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT0), .B(G128), .Z(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n194), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n257), .A2(new_n258), .A3(new_n253), .A4(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n244), .A2(new_n254), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(G110), .B(G140), .Z(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT79), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT70), .B(G953), .Z(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n272), .B(new_n274), .Z(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G469), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n257), .A2(new_n268), .A3(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n240), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n269), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n276), .A2(new_n277), .A3(new_n278), .A4(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n277), .A2(new_n278), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n270), .A2(new_n281), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n275), .A3(new_n269), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(G469), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT9), .B(G234), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT67), .B(G116), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G122), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n297), .A2(G122), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G107), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n201), .A3(new_n298), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT92), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT13), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n187), .A3(G128), .ZN(new_n305));
  XOR2_X1   g119(.A(G128), .B(G143), .Z(new_n306));
  OAI211_X1 g120(.A(G134), .B(new_n305), .C1(new_n306), .C2(new_n304), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n307), .A2(KEYINPUT93), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n306), .A2(G134), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n307), .B2(KEYINPUT93), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n300), .A2(new_n311), .A3(new_n301), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n303), .A2(new_n308), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n295), .A2(KEYINPUT14), .A3(G122), .ZN(new_n314));
  OAI211_X1 g128(.A(G107), .B(new_n314), .C1(new_n299), .C2(KEYINPUT14), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n306), .A2(G134), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n301), .C1(new_n309), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n291), .A2(new_n319), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n313), .A2(new_n317), .A3(new_n320), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n313), .A2(KEYINPUT94), .A3(new_n317), .A4(new_n320), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n278), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G478), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(KEYINPUT15), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n327), .A2(new_n328), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n332), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n339), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(G146), .ZN(new_n346));
  INV_X1    g160(.A(G237), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n273), .A2(G214), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(G143), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(new_n234), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT17), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n234), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n346), .B(new_n351), .C1(new_n352), .C2(KEYINPUT17), .ZN(new_n353));
  XNOR2_X1  g167(.A(G113), .B(G122), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(new_n204), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(KEYINPUT18), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT18), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n349), .B1(new_n357), .B2(new_n234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n342), .B(new_n190), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n345), .A2(new_n190), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n342), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n342), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(G146), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n362), .B(KEYINPUT91), .C1(G146), .C2(new_n366), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n352), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(new_n360), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n361), .B1(new_n372), .B2(new_n355), .ZN(new_n373));
  INV_X1    g187(.A(G475), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n278), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n361), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n355), .B1(new_n353), .B2(new_n360), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n278), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G475), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n373), .A2(KEYINPUT20), .A3(new_n374), .A4(new_n278), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n338), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  INV_X1    g199(.A(G952), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n386), .A2(KEYINPUT96), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(KEYINPUT96), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G234), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(new_n347), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT97), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n278), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT21), .B(G898), .Z(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G214), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  XOR2_X1   g215(.A(G110), .B(G122), .Z(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT8), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT67), .A2(G116), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT67), .A2(G116), .ZN(new_n405));
  OAI21_X1  g219(.A(G119), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n297), .A2(G119), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n408), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n297), .A2(KEYINPUT5), .A3(G119), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n410), .A2(KEYINPUT86), .ZN(new_n411));
  INV_X1    g225(.A(G113), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n410), .B2(KEYINPUT86), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n407), .B1(new_n295), .B2(G119), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT2), .B(G113), .Z(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n216), .A2(new_n418), .A3(KEYINPUT88), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT88), .B1(new_n216), .B2(new_n418), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n414), .A2(new_n417), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n218), .A2(new_n219), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n403), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n199), .A2(new_n339), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n385), .A2(G224), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n265), .A2(G125), .ZN(new_n427));
  AND4_X1   g241(.A1(KEYINPUT7), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n425), .A2(new_n427), .B1(KEYINPUT7), .B2(new_n426), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n401), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n221), .B2(new_n422), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n216), .A2(new_n418), .A3(KEYINPUT88), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n423), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n403), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n430), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT89), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n415), .B(new_n416), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n261), .A2(new_n440), .A3(new_n267), .ZN(new_n441));
  INV_X1    g255(.A(new_n402), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n423), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n431), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n423), .A2(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n402), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n425), .A2(new_n427), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(new_n426), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n445), .A2(new_n446), .A3(new_n451), .A4(new_n402), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n444), .A2(new_n453), .A3(new_n278), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n444), .A2(new_n453), .A3(new_n278), .A4(new_n455), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n398), .B(new_n400), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n294), .A2(new_n384), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n461));
  INV_X1    g275(.A(new_n199), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n227), .A2(KEYINPUT65), .A3(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n464), .C1(new_n229), .C2(G137), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G131), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n238), .B2(new_n239), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n251), .A2(new_n252), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT69), .A3(new_n466), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n473));
  INV_X1    g287(.A(new_n265), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n253), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n240), .A2(KEYINPUT68), .A3(new_n265), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n472), .A2(new_n477), .A3(new_n440), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT30), .B1(new_n472), .B2(new_n477), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n240), .A2(new_n265), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n199), .A3(new_n466), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n478), .B1(new_n484), .B2(new_n440), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n273), .A2(G210), .A3(new_n347), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT26), .B(G101), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n461), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n440), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n479), .B2(new_n483), .ZN(new_n494));
  NOR4_X1   g308(.A1(new_n494), .A2(KEYINPUT31), .A3(new_n490), .A4(new_n478), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n480), .B2(new_n482), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n478), .B2(new_n497), .ZN(new_n498));
  AOI221_X4 g312(.A(new_n468), .B1(new_n465), .B2(G131), .C1(new_n251), .C2(new_n252), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT69), .B1(new_n470), .B2(new_n466), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n199), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n493), .A3(new_n480), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n491), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n492), .A2(new_n495), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G472), .A2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT73), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n478), .ZN(new_n510));
  INV_X1    g324(.A(new_n483), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n475), .A3(new_n476), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(KEYINPUT30), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n491), .B(new_n510), .C1(new_n513), .C2(new_n493), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n498), .A2(new_n504), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n490), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n485), .A2(new_n461), .A3(new_n491), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT32), .B1(new_n519), .B2(new_n507), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n509), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n507), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n490), .B1(new_n494), .B2(new_n478), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(new_n516), .C2(new_n490), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n512), .A2(new_n440), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n510), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n491), .A2(KEYINPUT29), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n527), .B(new_n278), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n524), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT22), .Z(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n227), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G119), .ZN(new_n540));
  OR3_X1    g354(.A1(new_n540), .A2(KEYINPUT23), .A3(G128), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT23), .B1(new_n540), .B2(G128), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(new_n542), .B1(new_n540), .B2(G128), .ZN(new_n543));
  INV_X1    g357(.A(G110), .ZN(new_n544));
  XOR2_X1   g358(.A(G119), .B(G128), .Z(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT24), .B(G110), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n346), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n342), .A2(new_n190), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n550), .A2(new_n362), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n538), .A2(new_n548), .A3(new_n553), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n319), .B1(G234), .B2(new_n278), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G902), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT25), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n557), .A2(new_n278), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n278), .A3(new_n556), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n563), .B2(KEYINPUT25), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n558), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n460), .A2(new_n535), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(G101), .ZN(G3));
  INV_X1    g387(.A(new_n458), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n400), .B1(new_n574), .B2(KEYINPUT98), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n457), .A2(new_n576), .A3(new_n458), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n575), .B2(new_n577), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n325), .A2(new_n326), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n322), .A2(KEYINPUT33), .A3(new_n324), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G478), .A3(new_n278), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n327), .A2(new_n330), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n383), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n579), .A2(new_n580), .A3(new_n398), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n519), .B2(new_n278), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n523), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n593), .A2(new_n570), .A3(new_n293), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT34), .B(G104), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  INV_X1    g411(.A(new_n383), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n338), .ZN(new_n599));
  NOR4_X1   g413(.A1(new_n579), .A2(new_n580), .A3(new_n599), .A4(new_n398), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n594), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(new_n593), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n538), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT100), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n554), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n560), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n568), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n460), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT37), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n544), .ZN(G12));
  AND2_X1   g427(.A1(new_n609), .A2(new_n568), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n579), .A2(new_n580), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT101), .B(G900), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n394), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n393), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n615), .A2(new_n535), .A3(new_n294), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G128), .ZN(G30));
  NAND2_X1  g436(.A1(new_n457), .A2(new_n458), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT38), .Z(new_n624));
  NAND2_X1  g438(.A1(new_n338), .A2(new_n383), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n625), .A2(new_n610), .A3(new_n400), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n618), .B(KEYINPUT39), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n294), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT40), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n529), .A2(new_n490), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n514), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n632), .B2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n522), .A2(new_n524), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OR4_X1    g449(.A1(new_n624), .A2(new_n627), .A3(new_n630), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G143), .ZN(G45));
  NOR2_X1   g451(.A1(new_n588), .A2(new_n619), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n615), .A2(new_n535), .A3(new_n294), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G146), .ZN(G48));
  INV_X1    g454(.A(new_n589), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n276), .A2(new_n278), .A3(new_n282), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(G469), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(G469), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n276), .A2(new_n278), .A3(new_n282), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n292), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT104), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n644), .A2(new_n649), .A3(new_n292), .A4(new_n646), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n535), .A3(new_n571), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT105), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G15));
  NOR2_X1   g470(.A1(new_n579), .A2(new_n580), .ZN(new_n657));
  INV_X1    g471(.A(new_n398), .ZN(new_n658));
  INV_X1    g472(.A(new_n338), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n383), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n297), .ZN(G18));
  NOR3_X1   g477(.A1(new_n338), .A2(new_n383), .A3(new_n398), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n615), .A2(new_n651), .A3(new_n535), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT106), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n540), .ZN(G21));
  INV_X1    g481(.A(new_n625), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n492), .A2(new_n495), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n531), .A2(new_n490), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n508), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n591), .A2(new_n671), .A3(new_n570), .A4(new_n398), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n651), .A2(new_n657), .A3(new_n668), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G122), .ZN(G24));
  NOR2_X1   g488(.A1(new_n591), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n610), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n651), .A2(new_n677), .A3(new_n657), .A4(new_n638), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G125), .ZN(G27));
  NAND4_X1  g493(.A1(new_n280), .A2(KEYINPUT107), .A3(new_n275), .A4(new_n269), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n287), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n286), .A2(G469), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n283), .A3(new_n285), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n292), .A2(new_n399), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n457), .A2(new_n684), .A3(new_n458), .A4(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n535), .A2(new_n571), .A3(new_n638), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n638), .A2(new_n686), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n688), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT32), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n523), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n570), .B1(new_n695), .B2(new_n534), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n687), .A2(new_n688), .B1(new_n690), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n234), .ZN(G33));
  AND4_X1   g512(.A1(new_n535), .A2(new_n571), .A3(new_n620), .A4(new_n686), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n229), .ZN(G36));
  AOI21_X1  g514(.A(new_n383), .B1(new_n586), .B2(new_n585), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n383), .B2(KEYINPUT109), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n701), .B(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n593), .A3(new_n610), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n623), .A2(new_n400), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n288), .B1(new_n714), .B2(new_n277), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT108), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n286), .A2(KEYINPUT45), .A3(new_n680), .A4(new_n682), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n285), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n283), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(new_n292), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n712), .A2(new_n628), .A3(new_n713), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G137), .ZN(G39));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n292), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n638), .A2(new_n708), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n535), .A2(new_n730), .A3(new_n571), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(KEYINPUT111), .Z(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G140), .ZN(G42));
  INV_X1    g548(.A(new_n393), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n571), .A2(new_n704), .A3(new_n735), .A4(new_n675), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n644), .A2(new_n646), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n292), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n708), .B(new_n736), .C1(new_n729), .C2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n651), .A2(new_n708), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n571), .A3(new_n735), .A4(new_n635), .ZN(new_n741));
  OR3_X1    g555(.A1(new_n741), .A2(new_n383), .A3(new_n587), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n651), .A2(new_n400), .A3(new_n624), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT115), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n736), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n740), .A2(new_n735), .A3(new_n704), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n677), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n739), .A2(new_n742), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT51), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n665), .A2(new_n673), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n599), .A2(new_n588), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n594), .A2(new_n459), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n572), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n523), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n694), .B2(new_n509), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n570), .B1(new_n757), .B2(new_n534), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(new_n651), .C1(new_n600), .C2(new_n589), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n755), .A3(new_n759), .A4(new_n611), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n687), .A2(new_n688), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n690), .A2(new_n696), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n699), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n384), .A2(KEYINPUT113), .A3(new_n618), .A4(new_n708), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n535), .A2(new_n294), .A3(new_n610), .A4(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n338), .A2(new_n383), .A3(new_n619), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT113), .B1(new_n767), .B2(new_n708), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n689), .A2(new_n676), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n760), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n579), .A2(new_n580), .A3(new_n625), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n614), .A2(new_n618), .A3(new_n684), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n292), .A3(new_n634), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n621), .A2(new_n639), .A3(new_n775), .A4(new_n678), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n778), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n293), .B1(new_n757), .B2(new_n534), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(new_n615), .C1(new_n620), .C2(new_n638), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT52), .A3(new_n678), .A4(new_n775), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n783), .A3(KEYINPUT114), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n772), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n665), .A2(new_n673), .A3(new_n754), .A4(new_n572), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n652), .B1(new_n641), .B2(new_n661), .ZN(new_n789));
  INV_X1    g603(.A(new_n611), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n771), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n766), .A2(new_n768), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n697), .A2(new_n793), .A3(new_n699), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n780), .A2(new_n783), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n787), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n785), .A2(new_n786), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n779), .A3(new_n794), .A4(new_n792), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n780), .A2(new_n783), .A3(KEYINPUT114), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n787), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n780), .A2(new_n783), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n772), .A2(KEYINPUT53), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n786), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n748), .A2(new_n696), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n651), .A2(new_n657), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n389), .B1(new_n736), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n807), .B(new_n810), .C1(new_n588), .C2(new_n741), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT116), .Z(new_n812));
  NAND3_X1  g626(.A1(new_n751), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(G952), .B2(G953), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n737), .A2(KEYINPUT49), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n701), .A2(new_n816), .A3(new_n571), .A4(new_n685), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n634), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n815), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n737), .A2(KEYINPUT49), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n624), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(G75));
  AOI21_X1  g636(.A(new_n278), .B1(new_n785), .B2(new_n797), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(G210), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n450), .B(KEYINPUT55), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n448), .A2(new_n452), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT117), .Z(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n831), .B1(new_n829), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n273), .A2(G952), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G51));
  OR2_X1    g650(.A1(new_n285), .A2(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n285), .A2(KEYINPUT57), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n786), .B1(new_n785), .B2(new_n797), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n837), .B(new_n838), .C1(new_n798), .C2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n276), .A2(new_n282), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n840), .A2(KEYINPUT118), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n823), .A2(new_n717), .A3(new_n716), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(G54));
  NAND3_X1  g660(.A1(new_n823), .A2(KEYINPUT58), .A3(G475), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(new_n373), .Z(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n835), .ZN(G60));
  INV_X1    g663(.A(new_n584), .ZN(new_n850));
  NAND2_X1  g664(.A1(G478), .A2(G902), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT59), .Z(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n799), .A2(new_n800), .A3(new_n787), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT53), .B1(new_n772), .B2(new_n802), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n785), .A2(new_n797), .A3(new_n786), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT119), .B1(new_n859), .B2(new_n835), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n850), .B1(new_n805), .B2(new_n852), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n853), .B1(new_n798), .B2(new_n839), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n863));
  INV_X1    g677(.A(new_n835), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n860), .A2(new_n865), .A3(new_n861), .A4(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(G63));
  NAND2_X1  g684(.A1(G217), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT60), .Z(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n855), .B2(new_n856), .ZN(new_n873));
  INV_X1    g687(.A(new_n557), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n835), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n608), .B(KEYINPUT121), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g692(.A(new_n385), .B1(new_n395), .B2(G224), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n760), .B2(new_n273), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT122), .Z(new_n881));
  INV_X1    g695(.A(new_n831), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(G898), .B2(new_n273), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n881), .B(new_n883), .ZN(G69));
  XNOR2_X1  g698(.A(new_n484), .B(new_n366), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n724), .A2(new_n628), .A3(new_n696), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n887));
  INV_X1    g701(.A(new_n773), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n782), .A2(new_n678), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n763), .A3(new_n764), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n725), .A2(new_n733), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n273), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n895));
  XOR2_X1   g709(.A(KEYINPUT125), .B(G900), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n885), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n629), .A2(new_n623), .A3(new_n400), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n758), .A2(new_n753), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n636), .A2(new_n890), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n725), .A2(new_n733), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n636), .B(new_n890), .C1(KEYINPUT123), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n895), .B1(new_n908), .B2(new_n273), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n898), .B1(new_n909), .B2(new_n885), .ZN(G72));
  XNOR2_X1  g724(.A(new_n485), .B(KEYINPUT127), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n904), .A2(new_n760), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g726(.A1(G472), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT63), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT126), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n491), .B(new_n911), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n911), .A2(new_n491), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n891), .A2(new_n893), .A3(new_n760), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n801), .A2(new_n803), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n525), .A2(new_n514), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n864), .A2(new_n916), .A3(new_n919), .A4(new_n922), .ZN(G57));
endmodule


