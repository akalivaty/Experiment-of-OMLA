//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(G64gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT22), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n211), .A4(new_n214), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n208), .A2(new_n209), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n211), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT72), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT27), .B(G183gat), .Z(new_n225));
  OAI21_X1  g024(.A(KEYINPUT28), .B1(new_n225), .B2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  OR3_X1    g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT27), .B1(new_n227), .B2(new_n228), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n233), .A3(new_n234), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n231), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT24), .A3(new_n234), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n234), .A2(KEYINPUT24), .ZN(new_n249));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n243), .B(new_n247), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT65), .B(G169gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(KEYINPUT23), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(KEYINPUT23), .B1(new_n236), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n249), .A2(new_n250), .ZN(new_n259));
  INV_X1    g058(.A(new_n247), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n256), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n235), .B2(KEYINPUT23), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n261), .A2(KEYINPUT66), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n262), .A2(new_n245), .A3(new_n247), .A4(new_n264), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n242), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT73), .B(new_n242), .C1(new_n258), .C2(new_n269), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT74), .ZN(new_n278));
  INV_X1    g077(.A(new_n242), .ZN(new_n279));
  INV_X1    g078(.A(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n255), .A2(KEYINPUT23), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT64), .B1(new_n259), .B2(new_n260), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n262), .A4(new_n251), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n263), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n279), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n285), .B2(new_n276), .ZN(new_n286));
  INV_X1    g085(.A(new_n276), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n224), .B1(new_n277), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n222), .B(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n274), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n285), .A2(KEYINPUT29), .A3(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n207), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n276), .B1(new_n272), .B2(new_n274), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n224), .B1(new_n298), .B2(new_n294), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n275), .A2(new_n276), .B1(new_n286), .B2(new_n288), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n299), .B(new_n206), .C1(new_n300), .C2(new_n224), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(KEYINPUT30), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(new_n300), .B2(new_n224), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n207), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(KEYINPUT82), .A3(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n321), .A2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n316), .A2(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n317), .A2(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n323), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G113gat), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n341), .A2(new_n339), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT69), .A3(new_n338), .A4(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT1), .B1(new_n334), .B2(new_n336), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n324), .A2(new_n328), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n332), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT70), .B1(new_n347), .B2(new_n350), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n360), .B(new_n349), .C1(new_n344), .C2(new_n346), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n358), .B(new_n353), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n353), .A2(new_n347), .A3(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n362), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT78), .B1(new_n362), .B2(new_n364), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n354), .B(new_n357), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n347), .A2(KEYINPUT70), .A3(new_n350), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n356), .B1(new_n363), .B2(new_n358), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n354), .ZN(new_n373));
  INV_X1    g172(.A(new_n353), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n363), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n356), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(KEYINPUT5), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n311), .B1(new_n367), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT83), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n378), .A3(new_n311), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT39), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n356), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n354), .B1(new_n365), .B2(new_n366), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n356), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n391), .A3(new_n356), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n386), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT40), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n390), .B(KEYINPUT40), .C1(new_n394), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n310), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n277), .A2(new_n289), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n224), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n291), .B1(new_n298), .B2(new_n294), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT86), .B(new_n291), .C1(new_n298), .C2(new_n294), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT37), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n303), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT38), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(KEYINPUT87), .A3(KEYINPUT37), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n206), .A4(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n297), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n207), .B1(new_n303), .B2(new_n411), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n299), .B(KEYINPUT37), .C1(new_n300), .C2(new_n224), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n412), .A2(new_n420), .A3(new_n206), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT38), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT88), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n367), .A2(new_n378), .ZN(new_n428));
  INV_X1    g227(.A(new_n385), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n385), .B1(new_n367), .B2(new_n378), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n389), .A2(new_n431), .B1(KEYINPUT6), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n423), .A3(new_n426), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n219), .A2(new_n221), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT79), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n215), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n273), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n353), .B1(new_n440), .B2(new_n331), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n332), .A2(new_n273), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n224), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G228gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n352), .B1(new_n222), .B2(KEYINPUT29), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n449), .B2(new_n374), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n332), .A2(KEYINPUT80), .A3(new_n273), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n324), .A2(new_n328), .A3(new_n330), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(KEYINPUT29), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n450), .B1(new_n455), .B2(new_n291), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n443), .B2(new_n445), .ZN(new_n458));
  OAI21_X1  g257(.A(G22gat), .B1(new_n458), .B2(KEYINPUT81), .ZN(new_n459));
  XOR2_X1   g258(.A(G78gat), .B(G106gat), .Z(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n458), .B2(KEYINPUT81), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n457), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n459), .B2(new_n457), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n402), .A2(new_n434), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n430), .B(new_n432), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n306), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n370), .A2(new_n270), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n359), .A2(new_n361), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n285), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  INV_X1    g274(.A(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT34), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT32), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n474), .ZN(new_n483));
  INV_X1    g282(.A(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n480), .B2(new_n482), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G71gat), .ZN(new_n489));
  INV_X1    g288(.A(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n478), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(KEYINPUT33), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n486), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  INV_X1    g294(.A(new_n482), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n481), .B1(new_n478), .B2(KEYINPUT32), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n484), .B(new_n483), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT36), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n494), .B2(new_n500), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n469), .A2(new_n471), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n468), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g307(.A(new_n388), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n509), .A2(new_n379), .A3(new_n386), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n510), .B2(new_n430), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n308), .A3(new_n309), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n493), .B1(new_n486), .B2(new_n487), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n495), .A3(new_n499), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n467), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n507), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n467), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT35), .B1(new_n471), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n302), .A2(KEYINPUT82), .A3(new_n305), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT82), .B1(new_n302), .B2(new_n305), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT89), .A4(new_n511), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n527), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT93), .B(G8gat), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n534), .B1(new_n530), .B2(new_n531), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT94), .A3(new_n533), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n530), .A2(G8gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT14), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n554));
  INV_X1    g353(.A(new_n544), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n538), .A2(new_n540), .B1(G8gat), .B2(new_n530), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n553), .A2(new_n562), .A3(new_n556), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT18), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n557), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n565), .B(KEYINPUT13), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT91), .B(G169gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n583), .A3(new_n573), .A4(new_n575), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n526), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G64gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G78gat), .ZN(new_n593));
  AND2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n593), .ZN(new_n597));
  OR2_X1    g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT9), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(KEYINPUT98), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT20), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n560), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n616), .A2(KEYINPUT100), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT19), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(KEYINPUT100), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT19), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(KEYINPUT20), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT99), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n622), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n622), .B2(new_n626), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n613), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n622), .A2(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n628), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n622), .A2(new_n626), .A3(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n612), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(G99gat), .A2(G106gat), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n640), .B1(new_n641), .B2(new_n205), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G99gat), .B(G106gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n642), .A3(new_n639), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n561), .A2(new_n648), .A3(new_n563), .ZN(new_n649));
  NAND3_X1  g448(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n645), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n558), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G190gat), .B(G218gat), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n653), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT102), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n649), .A2(new_n652), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n661), .A2(KEYINPUT101), .A3(new_n650), .A4(new_n655), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT102), .B(new_n670), .C1(new_n658), .C2(new_n659), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n637), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  INV_X1    g475(.A(new_n602), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n651), .A2(KEYINPUT104), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n648), .B2(new_n602), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n606), .B2(new_n648), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n596), .A2(KEYINPUT98), .A3(new_n601), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n596), .B2(new_n601), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n682), .B(new_n648), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n676), .B(new_n681), .C1(new_n683), .C2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n651), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n675), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n681), .B1(new_n683), .B2(new_n687), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n675), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT106), .ZN(new_n696));
  INV_X1    g495(.A(G176gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(G204gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n526), .A2(KEYINPUT96), .A3(new_n587), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n590), .A2(new_n673), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n470), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g511(.A(G8gat), .B1(new_n708), .B2(new_n523), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT96), .B1(new_n526), .B2(new_n587), .ZN(new_n714));
  INV_X1    g513(.A(new_n587), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n589), .B(new_n715), .C1(new_n506), .C2(new_n525), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n714), .A2(new_n716), .A3(new_n705), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT107), .B(G8gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n528), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n673), .A3(new_n310), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n713), .B2(new_n720), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n523), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT42), .B1(new_n728), .B2(new_n719), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT108), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1325gat));
  INV_X1    g530(.A(G15gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n502), .A2(new_n504), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n708), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n709), .A2(new_n501), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n732), .ZN(G1326gat));
  NOR2_X1   g535(.A1(new_n708), .A2(new_n467), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT43), .B(G22gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1327gat));
  INV_X1    g538(.A(new_n672), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n714), .A2(new_n716), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n637), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n705), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(G29gat), .A3(new_n470), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n746));
  OR2_X1    g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n526), .A2(new_n672), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n526), .A2(new_n751), .A3(KEYINPUT44), .A4(new_n672), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n750), .A2(new_n587), .A3(new_n743), .A4(new_n752), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n753), .A2(KEYINPUT111), .A3(new_n470), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT111), .B1(new_n753), .B2(new_n470), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(G29gat), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n745), .A2(new_n746), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n747), .A2(new_n756), .A3(new_n757), .ZN(G1328gat));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n546), .A3(new_n310), .A4(new_n743), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n753), .B2(new_n523), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(G1329gat));
  OAI21_X1  g562(.A(G43gat), .B1(new_n753), .B2(new_n733), .ZN(new_n764));
  INV_X1    g563(.A(G43gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n741), .A2(new_n765), .A3(new_n501), .A4(new_n743), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g567(.A(G50gat), .B1(new_n753), .B2(new_n467), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT48), .B1(new_n769), .B2(KEYINPUT112), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n467), .A2(G50gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n744), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n770), .B(new_n772), .ZN(G1331gat));
  NAND3_X1  g572(.A1(new_n673), .A2(new_n705), .A3(new_n715), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n673), .A2(KEYINPUT113), .A3(new_n705), .A4(new_n715), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n776), .A2(new_n777), .B1(new_n506), .B2(new_n525), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n710), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n778), .B(new_n310), .C1(new_n781), .C2(new_n203), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT114), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n203), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1333gat));
  INV_X1    g584(.A(new_n733), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n778), .A2(G71gat), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n778), .A2(new_n501), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(G71gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n778), .A2(new_n469), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n742), .A2(new_n587), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n526), .A2(new_n672), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n706), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n641), .A3(new_n710), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n750), .A2(new_n705), .A3(new_n752), .A4(new_n793), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n470), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1336gat));
  OAI21_X1  g601(.A(G92gat), .B1(new_n800), .B2(new_n523), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n795), .B2(new_n796), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n794), .A2(KEYINPUT116), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n310), .A2(new_n205), .A3(new_n705), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(KEYINPUT115), .B(G92gat), .C1(new_n800), .C2(new_n523), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n805), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n816));
  OAI211_X1 g615(.A(new_n803), .B(new_n816), .C1(new_n797), .C2(new_n810), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1337gat));
  NOR3_X1   g617(.A1(new_n800), .A2(new_n490), .A3(new_n733), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n501), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n490), .ZN(G1338gat));
  NOR3_X1   g620(.A1(new_n706), .A2(G106gat), .A3(new_n467), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n807), .A2(new_n809), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n800), .A2(new_n467), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  INV_X1    g627(.A(new_n822), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n797), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n826), .B2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n688), .A2(new_n675), .A3(new_n689), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n690), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n690), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n838), .B2(new_n701), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT118), .B(new_n700), .C1(new_n690), .C2(new_n837), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT54), .B(new_n675), .C1(new_n688), .C2(new_n689), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n844), .B2(new_n700), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n836), .A3(new_n701), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT55), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n843), .A2(new_n703), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n571), .A2(new_n572), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n565), .B1(new_n559), .B2(new_n564), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n582), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n586), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n849), .A2(KEYINPUT119), .A3(new_n672), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n702), .B1(new_n847), .B2(KEYINPUT55), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n672), .A2(new_n855), .A3(new_n853), .A4(new_n843), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n705), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n843), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n715), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n740), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n742), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NOR4_X1   g663(.A1(new_n637), .A2(new_n672), .A3(new_n705), .A4(new_n587), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n310), .A2(new_n470), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n866), .A2(new_n518), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n587), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n705), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n742), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(G127gat), .ZN(G1342gat));
  NOR3_X1   g674(.A1(new_n866), .A2(new_n740), .A3(new_n868), .ZN(new_n876));
  INV_X1    g675(.A(new_n518), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT56), .B(G134gat), .Z(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n841), .A2(KEYINPUT121), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n847), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n884), .A3(new_n842), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n587), .A3(new_n855), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n860), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n740), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n742), .B1(new_n888), .B2(new_n859), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT57), .B(new_n469), .C1(new_n889), .C2(new_n865), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT122), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n866), .B2(new_n467), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n673), .A2(new_n706), .A3(new_n715), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n740), .A2(new_n887), .B1(new_n854), .B2(new_n858), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n742), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT57), .A4(new_n469), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n868), .A2(new_n786), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n587), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n866), .A2(new_n467), .A3(new_n786), .A4(new_n868), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n313), .A3(new_n587), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  OAI211_X1 g709(.A(new_n469), .B(new_n892), .C1(new_n864), .C2(new_n865), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n672), .B1(new_n886), .B2(new_n860), .ZN(new_n912));
  INV_X1    g711(.A(new_n856), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n637), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n467), .B1(new_n914), .B2(new_n895), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(KEYINPUT57), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n705), .A3(new_n901), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n904), .B2(new_n705), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n901), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n705), .A2(new_n919), .ZN(new_n922));
  OAI221_X1 g721(.A(new_n918), .B1(new_n920), .B2(G148gat), .C1(new_n921), .C2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n921), .B2(new_n637), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n319), .A3(new_n742), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(KEYINPUT123), .B1(new_n921), .B2(new_n740), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n900), .A2(new_n928), .A3(new_n672), .A4(new_n901), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(G162gat), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n876), .A2(new_n320), .A3(new_n469), .A4(new_n733), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n866), .A2(new_n710), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n310), .A3(new_n877), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  INV_X1    g734(.A(new_n254), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n587), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n934), .B2(new_n715), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n934), .A2(new_n697), .A3(new_n706), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n935), .A2(new_n705), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n697), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n934), .A2(new_n637), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n225), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n228), .B1(new_n934), .B2(new_n637), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n934), .B2(new_n740), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n231), .A3(new_n672), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n733), .A2(new_n310), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(new_n710), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n916), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n715), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n953), .B2(new_n467), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n733), .A2(KEYINPUT125), .A3(new_n469), .A4(new_n310), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n933), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n715), .A2(G197gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  NOR3_X1   g762(.A1(new_n961), .A2(G204gat), .A3(new_n706), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g766(.A(G204gat), .B1(new_n956), .B2(new_n706), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n916), .A2(new_n742), .A3(new_n954), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n916), .A2(new_n972), .A3(new_n742), .A4(new_n954), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(G211gat), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n961), .A2(G211gat), .A3(new_n637), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1354gat));
  NOR3_X1   g779(.A1(new_n956), .A2(new_n213), .A3(new_n740), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n961), .A2(new_n740), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n213), .B2(new_n982), .ZN(G1355gat));
endmodule


