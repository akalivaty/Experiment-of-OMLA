

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781;

  NAND2_X1 U370 ( .A1(n348), .A2(n669), .ZN(n672) );
  AND2_X1 U371 ( .A1(n377), .A2(n535), .ZN(n376) );
  NOR2_X1 U372 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U373 ( .A(n546), .ZN(n554) );
  NAND2_X1 U374 ( .A1(n424), .A2(n365), .ZN(n411) );
  XNOR2_X1 U375 ( .A(n520), .B(KEYINPUT97), .ZN(n768) );
  XNOR2_X1 U376 ( .A(n423), .B(n422), .ZN(n763) );
  XNOR2_X1 U377 ( .A(n428), .B(n427), .ZN(n769) );
  NAND2_X2 U378 ( .A1(n350), .A2(n351), .ZN(n551) );
  AND2_X1 U379 ( .A1(n347), .A2(n720), .ZN(n557) );
  XNOR2_X1 U380 ( .A(n388), .B(KEYINPUT108), .ZN(n347) );
  NAND2_X1 U381 ( .A1(n668), .A2(n667), .ZN(n348) );
  XNOR2_X1 U382 ( .A(n769), .B(G146), .ZN(n491) );
  NAND2_X1 U383 ( .A1(n673), .A2(n674), .ZN(n584) );
  INV_X1 U384 ( .A(n584), .ZN(n676) );
  AND2_X2 U385 ( .A1(n634), .A2(n669), .ZN(n749) );
  BUF_X1 U386 ( .A(n749), .Z(n349) );
  INV_X1 U387 ( .A(G953), .ZN(n771) );
  NAND2_X2 U388 ( .A1(n352), .A2(n353), .ZN(n393) );
  NAND2_X1 U389 ( .A1(n542), .A2(n544), .ZN(n600) );
  NOR2_X2 U390 ( .A1(G953), .A2(G237), .ZN(n510) );
  XNOR2_X1 U391 ( .A(n682), .B(KEYINPUT6), .ZN(n615) );
  XNOR2_X1 U392 ( .A(n482), .B(n389), .ZN(n544) );
  XNOR2_X1 U393 ( .A(n518), .B(G472), .ZN(n682) );
  XNOR2_X1 U394 ( .A(n768), .B(n526), .ZN(n745) );
  XNOR2_X1 U395 ( .A(n447), .B(G146), .ZN(n508) );
  XNOR2_X1 U396 ( .A(n452), .B(n513), .ZN(n525) );
  INV_X2 U397 ( .A(KEYINPUT3), .ZN(n410) );
  INV_X1 U398 ( .A(KEYINPUT4), .ZN(n447) );
  XNOR2_X1 U399 ( .A(G128), .B(G137), .ZN(n494) );
  XNOR2_X2 U400 ( .A(KEYINPUT10), .B(G140), .ZN(n428) );
  AND2_X1 U401 ( .A1(n373), .A2(n372), .ZN(n350) );
  OR2_X1 U402 ( .A1(n745), .A2(n369), .ZN(n351) );
  NAND2_X1 U403 ( .A1(n404), .A2(KEYINPUT34), .ZN(n352) );
  AND2_X1 U404 ( .A1(n354), .A2(n405), .ZN(n353) );
  INV_X1 U405 ( .A(n394), .ZN(n354) );
  AND2_X2 U406 ( .A1(n617), .A2(n437), .ZN(n417) );
  AND2_X1 U407 ( .A1(n416), .A2(n533), .ZN(n363) );
  AND2_X2 U408 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X2 U409 ( .A(n506), .B(n434), .ZN(n673) );
  NOR2_X1 U410 ( .A1(n660), .A2(n664), .ZN(n633) );
  INV_X1 U411 ( .A(n598), .ZN(n688) );
  XNOR2_X1 U412 ( .A(n383), .B(n382), .ZN(n562) );
  INV_X1 U413 ( .A(KEYINPUT71), .ZN(n382) );
  XOR2_X1 U414 ( .A(G107), .B(G122), .Z(n469) );
  XOR2_X1 U415 ( .A(G104), .B(G113), .Z(n473) );
  XNOR2_X1 U416 ( .A(G902), .B(KEYINPUT15), .ZN(n629) );
  XNOR2_X1 U417 ( .A(G137), .B(G131), .ZN(n507) );
  AND2_X1 U418 ( .A1(n598), .A2(n613), .ZN(n599) );
  AND2_X1 U419 ( .A1(n689), .A2(n674), .ZN(n380) );
  NAND2_X1 U420 ( .A1(n465), .A2(n357), .ZN(n425) );
  XNOR2_X1 U421 ( .A(n468), .B(n442), .ZN(n441) );
  INV_X1 U422 ( .A(KEYINPUT7), .ZN(n442) );
  XNOR2_X1 U423 ( .A(KEYINPUT70), .B(G110), .ZN(n452) );
  XNOR2_X1 U424 ( .A(n431), .B(n367), .ZN(n623) );
  XNOR2_X1 U425 ( .A(n438), .B(n358), .ZN(n542) );
  XNOR2_X1 U426 ( .A(n653), .B(n652), .ZN(n654) );
  AND2_X1 U427 ( .A1(n781), .A2(n355), .ZN(n381) );
  AND2_X1 U428 ( .A1(n781), .A2(n726), .ZN(n537) );
  INV_X1 U429 ( .A(KEYINPUT89), .ZN(n407) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n458) );
  OR2_X1 U431 ( .A1(G902), .A2(G237), .ZN(n455) );
  NAND2_X1 U432 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U433 ( .A(n527), .ZN(n371) );
  XNOR2_X1 U434 ( .A(KEYINPUT5), .B(G113), .ZN(n511) );
  INV_X1 U435 ( .A(G125), .ZN(n427) );
  XOR2_X1 U436 ( .A(KEYINPUT103), .B(G122), .Z(n478) );
  XNOR2_X1 U437 ( .A(G143), .B(G131), .ZN(n477) );
  XOR2_X1 U438 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n475) );
  NOR2_X1 U439 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U440 ( .A(G125), .B(KEYINPUT17), .ZN(n450) );
  XNOR2_X1 U441 ( .A(n508), .B(n448), .ZN(n449) );
  NAND2_X1 U442 ( .A1(n386), .A2(n391), .ZN(n415) );
  AND2_X1 U443 ( .A1(n356), .A2(n436), .ZN(n386) );
  INV_X1 U444 ( .A(KEYINPUT38), .ZN(n387) );
  INV_X1 U445 ( .A(KEYINPUT19), .ZN(n457) );
  OR2_X1 U446 ( .A1(n635), .A2(G902), .ZN(n518) );
  XNOR2_X1 U447 ( .A(n564), .B(KEYINPUT45), .ZN(n565) );
  XNOR2_X1 U448 ( .A(n453), .B(n473), .ZN(n422) );
  XNOR2_X1 U449 ( .A(n515), .B(n454), .ZN(n423) );
  XNOR2_X1 U450 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U451 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U452 ( .A(KEYINPUT24), .ZN(n496) );
  XNOR2_X1 U453 ( .A(KEYINPUT100), .B(KEYINPUT23), .ZN(n492) );
  XOR2_X1 U454 ( .A(KEYINPUT98), .B(KEYINPUT74), .Z(n493) );
  XNOR2_X1 U455 ( .A(n763), .B(n418), .ZN(n644) );
  XNOR2_X1 U456 ( .A(n421), .B(n419), .ZN(n418) );
  XNOR2_X1 U457 ( .A(n449), .B(n525), .ZN(n421) );
  XNOR2_X1 U458 ( .A(n420), .B(n451), .ZN(n419) );
  NAND2_X1 U459 ( .A1(n582), .A2(n613), .ZN(n406) );
  AND2_X1 U460 ( .A1(n588), .A2(n432), .ZN(n594) );
  INV_X1 U461 ( .A(n589), .ZN(n433) );
  BUF_X1 U462 ( .A(n682), .Z(n385) );
  XNOR2_X1 U463 ( .A(n483), .B(n484), .ZN(n389) );
  INV_X1 U464 ( .A(KEYINPUT22), .ZN(n488) );
  AND2_X1 U465 ( .A1(n411), .A2(n380), .ZN(n379) );
  BUF_X1 U466 ( .A(n391), .Z(n390) );
  XNOR2_X1 U467 ( .A(n505), .B(KEYINPUT25), .ZN(n434) );
  XNOR2_X1 U468 ( .A(n635), .B(KEYINPUT62), .ZN(n636) );
  XNOR2_X1 U469 ( .A(n443), .B(n440), .ZN(n472) );
  XNOR2_X1 U470 ( .A(n470), .B(n441), .ZN(n440) );
  NAND2_X1 U471 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U472 ( .A(G140), .B(G107), .ZN(n522) );
  AND2_X1 U473 ( .A1(n638), .A2(G953), .ZN(n753) );
  AND2_X1 U474 ( .A1(n726), .A2(n368), .ZN(n355) );
  XNOR2_X1 U475 ( .A(n406), .B(n457), .ZN(n575) );
  AND2_X1 U476 ( .A1(n676), .A2(KEYINPUT33), .ZN(n356) );
  XOR2_X1 U477 ( .A(n466), .B(KEYINPUT0), .Z(n357) );
  XOR2_X1 U478 ( .A(KEYINPUT106), .B(G478), .Z(n358) );
  XOR2_X1 U479 ( .A(n508), .B(n507), .Z(n359) );
  BUF_X1 U480 ( .A(n661), .Z(n754) );
  AND2_X1 U481 ( .A1(n435), .A2(n437), .ZN(n360) );
  XOR2_X1 U482 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n361) );
  OR2_X1 U483 ( .A1(n612), .A2(n406), .ZN(n362) );
  INV_X1 U484 ( .A(n674), .ZN(n439) );
  NAND2_X1 U485 ( .A1(n412), .A2(n411), .ZN(n546) );
  AND2_X1 U486 ( .A1(n591), .A2(n398), .ZN(n364) );
  NOR2_X1 U487 ( .A1(n465), .A2(n357), .ZN(n365) );
  NOR2_X1 U488 ( .A1(n673), .A2(n385), .ZN(n366) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(n595), .Z(n367) );
  INV_X1 U490 ( .A(G902), .ZN(n370) );
  INV_X1 U491 ( .A(KEYINPUT33), .ZN(n437) );
  AND2_X1 U492 ( .A1(n536), .A2(KEYINPUT44), .ZN(n368) );
  XNOR2_X2 U493 ( .A(n551), .B(n392), .ZN(n617) );
  NAND2_X1 U494 ( .A1(n527), .A2(G902), .ZN(n372) );
  NAND2_X1 U495 ( .A1(n745), .A2(n527), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n376), .A2(n374), .ZN(n558) );
  NAND2_X1 U497 ( .A1(n375), .A2(n537), .ZN(n374) );
  NOR2_X1 U498 ( .A1(n715), .A2(n536), .ZN(n375) );
  NAND2_X1 U499 ( .A1(n381), .A2(n715), .ZN(n377) );
  XNOR2_X2 U500 ( .A(n378), .B(n488), .ZN(n540) );
  NAND2_X1 U501 ( .A1(n379), .A2(n412), .ZN(n378) );
  NAND2_X1 U502 ( .A1(n402), .A2(n534), .ZN(n397) );
  NAND2_X1 U503 ( .A1(n403), .A2(n405), .ZN(n402) );
  XNOR2_X1 U504 ( .A(n559), .B(KEYINPUT87), .ZN(n563) );
  NAND2_X1 U505 ( .A1(n561), .A2(n560), .ZN(n383) );
  XNOR2_X2 U506 ( .A(n384), .B(n565), .ZN(n661) );
  NAND2_X1 U507 ( .A1(n563), .A2(n562), .ZN(n384) );
  AND2_X2 U508 ( .A1(n426), .A2(n425), .ZN(n412) );
  XNOR2_X2 U509 ( .A(n621), .B(n387), .ZN(n598) );
  NAND2_X1 U510 ( .A1(n555), .A2(n576), .ZN(n388) );
  XNOR2_X1 U511 ( .A(n479), .B(n445), .ZN(n480) );
  XNOR2_X1 U512 ( .A(n481), .B(n480), .ZN(n653) );
  NAND2_X1 U513 ( .A1(n633), .A2(n430), .ZN(n669) );
  INV_X1 U514 ( .A(n617), .ZN(n391) );
  OR2_X1 U515 ( .A1(n617), .A2(n584), .ZN(n547) );
  AND2_X1 U516 ( .A1(n617), .A2(n366), .ZN(n532) );
  AND2_X1 U517 ( .A1(n617), .A2(n584), .ZN(n677) );
  NOR2_X1 U518 ( .A1(n390), .A2(n538), .ZN(n539) );
  AND2_X1 U519 ( .A1(n580), .A2(n390), .ZN(n739) );
  INV_X1 U520 ( .A(KEYINPUT1), .ZN(n392) );
  NAND2_X2 U521 ( .A1(n395), .A2(n393), .ZN(n715) );
  NAND2_X1 U522 ( .A1(n400), .A2(n364), .ZN(n394) );
  NAND2_X1 U523 ( .A1(n399), .A2(n534), .ZN(n396) );
  INV_X1 U524 ( .A(n414), .ZN(n404) );
  INV_X1 U525 ( .A(n534), .ZN(n398) );
  NAND2_X1 U526 ( .A1(n400), .A2(n591), .ZN(n399) );
  NAND2_X1 U527 ( .A1(n401), .A2(KEYINPUT34), .ZN(n400) );
  INV_X1 U528 ( .A(n416), .ZN(n401) );
  NAND2_X1 U529 ( .A1(n404), .A2(KEYINPUT34), .ZN(n403) );
  NAND2_X1 U530 ( .A1(n363), .A2(n414), .ZN(n405) );
  XNOR2_X1 U531 ( .A(n537), .B(n407), .ZN(n561) );
  XNOR2_X2 U532 ( .A(n409), .B(n408), .ZN(n515) );
  XNOR2_X2 U533 ( .A(G119), .B(G116), .ZN(n408) );
  XNOR2_X2 U534 ( .A(n410), .B(KEYINPUT69), .ZN(n409) );
  XNOR2_X2 U535 ( .A(n413), .B(G143), .ZN(n471) );
  XNOR2_X2 U536 ( .A(G128), .B(KEYINPUT77), .ZN(n413) );
  NAND2_X1 U537 ( .A1(n416), .A2(n415), .ZN(n705) );
  AND2_X2 U538 ( .A1(n415), .A2(n554), .ZN(n414) );
  NOR2_X2 U539 ( .A1(n360), .A2(n417), .ZN(n416) );
  INV_X1 U540 ( .A(n471), .ZN(n420) );
  INV_X1 U541 ( .A(n575), .ZN(n424) );
  NAND2_X1 U542 ( .A1(n575), .A2(n357), .ZN(n426) );
  XNOR2_X2 U543 ( .A(KEYINPUT67), .B(G101), .ZN(n513) );
  INV_X1 U544 ( .A(n770), .ZN(n660) );
  NAND2_X1 U545 ( .A1(n429), .A2(n664), .ZN(n663) );
  NAND2_X1 U546 ( .A1(n430), .A2(n770), .ZN(n429) );
  INV_X1 U547 ( .A(n661), .ZN(n430) );
  NAND2_X1 U548 ( .A1(n594), .A2(n598), .ZN(n431) );
  AND2_X1 U549 ( .A1(n587), .A2(n433), .ZN(n432) );
  XNOR2_X2 U550 ( .A(n509), .B(n359), .ZN(n520) );
  XNOR2_X2 U551 ( .A(n471), .B(G134), .ZN(n509) );
  NAND2_X1 U552 ( .A1(n436), .A2(n676), .ZN(n435) );
  INV_X1 U553 ( .A(n615), .ZN(n436) );
  INV_X1 U554 ( .A(n542), .ZN(n545) );
  NAND2_X1 U555 ( .A1(n751), .A2(n370), .ZN(n438) );
  NAND2_X1 U556 ( .A1(n540), .A2(n530), .ZN(n531) );
  NAND2_X1 U557 ( .A1(n489), .A2(G217), .ZN(n443) );
  AND2_X1 U558 ( .A1(G210), .A2(n455), .ZN(n444) );
  XOR2_X1 U559 ( .A(n478), .B(n477), .Z(n445) );
  XNOR2_X1 U560 ( .A(n608), .B(KEYINPUT46), .ZN(n609) );
  INV_X1 U561 ( .A(n469), .ZN(n454) );
  NAND2_X1 U562 ( .A1(G214), .A2(n455), .ZN(n446) );
  XNOR2_X1 U563 ( .A(KEYINPUT92), .B(n446), .ZN(n613) );
  NAND2_X1 U564 ( .A1(G224), .A2(n771), .ZN(n448) );
  XNOR2_X1 U565 ( .A(n361), .B(n450), .ZN(n451) );
  XOR2_X1 U566 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n453) );
  NAND2_X1 U567 ( .A1(n644), .A2(n629), .ZN(n456) );
  XNOR2_X2 U568 ( .A(n456), .B(n444), .ZN(n582) );
  XNOR2_X1 U569 ( .A(n458), .B(KEYINPUT14), .ZN(n459) );
  NAND2_X1 U570 ( .A1(n459), .A2(G952), .ZN(n702) );
  NOR2_X1 U571 ( .A1(G953), .A2(n702), .ZN(n569) );
  XOR2_X1 U572 ( .A(KEYINPUT93), .B(G898), .Z(n761) );
  NAND2_X1 U573 ( .A1(G902), .A2(n459), .ZN(n460) );
  XOR2_X1 U574 ( .A(KEYINPUT94), .B(n460), .Z(n461) );
  NAND2_X1 U575 ( .A1(G953), .A2(n461), .ZN(n567) );
  NOR2_X1 U576 ( .A1(n761), .A2(n567), .ZN(n462) );
  XOR2_X1 U577 ( .A(KEYINPUT95), .B(n462), .Z(n463) );
  NOR2_X1 U578 ( .A1(n569), .A2(n463), .ZN(n464) );
  XNOR2_X1 U579 ( .A(n464), .B(KEYINPUT96), .ZN(n465) );
  INV_X1 U580 ( .A(KEYINPUT90), .ZN(n466) );
  XOR2_X1 U581 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n468) );
  NAND2_X1 U582 ( .A1(G234), .A2(n771), .ZN(n467) );
  XOR2_X1 U583 ( .A(KEYINPUT8), .B(n467), .Z(n489) );
  XNOR2_X1 U584 ( .A(G116), .B(n469), .ZN(n470) );
  XNOR2_X1 U585 ( .A(n509), .B(n472), .ZN(n751) );
  XNOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n491), .B(n473), .ZN(n481) );
  NAND2_X1 U588 ( .A1(G214), .A2(n510), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U590 ( .A(n476), .B(KEYINPUT12), .Z(n479) );
  NOR2_X1 U591 ( .A1(G902), .A2(n653), .ZN(n482) );
  INV_X1 U592 ( .A(G475), .ZN(n484) );
  INV_X1 U593 ( .A(n600), .ZN(n689) );
  NAND2_X1 U594 ( .A1(n629), .A2(G234), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n485), .B(KEYINPUT20), .ZN(n504) );
  NAND2_X1 U596 ( .A1(n504), .A2(G221), .ZN(n487) );
  INV_X1 U597 ( .A(KEYINPUT21), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n487), .B(n486), .ZN(n674) );
  NAND2_X1 U599 ( .A1(G221), .A2(n489), .ZN(n490) );
  XNOR2_X1 U600 ( .A(n491), .B(n490), .ZN(n503) );
  XOR2_X1 U601 ( .A(n493), .B(n492), .Z(n501) );
  XOR2_X1 U602 ( .A(KEYINPUT80), .B(KEYINPUT99), .Z(n495) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n499) );
  XNOR2_X1 U604 ( .A(G110), .B(G119), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U606 ( .A(n502), .B(n503), .ZN(n716) );
  NOR2_X1 U607 ( .A1(G902), .A2(n716), .ZN(n506) );
  NAND2_X1 U608 ( .A1(G217), .A2(n504), .ZN(n505) );
  INV_X1 U609 ( .A(n673), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n510), .A2(G210), .ZN(n512) );
  XNOR2_X1 U611 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n515), .B(n516), .ZN(n517) );
  XNOR2_X1 U614 ( .A(n520), .B(n517), .ZN(n635) );
  NAND2_X1 U615 ( .A1(n519), .A2(n615), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n771), .A2(G227), .ZN(n521) );
  XNOR2_X1 U617 ( .A(n521), .B(G104), .ZN(n523) );
  XNOR2_X1 U618 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U619 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U620 ( .A(KEYINPUT68), .B(G469), .ZN(n527) );
  NOR2_X1 U621 ( .A1(n528), .A2(n617), .ZN(n529) );
  XNOR2_X1 U622 ( .A(n529), .B(KEYINPUT76), .ZN(n530) );
  XNOR2_X2 U623 ( .A(n531), .B(KEYINPUT32), .ZN(n781) );
  NAND2_X1 U624 ( .A1(n540), .A2(n532), .ZN(n726) );
  INV_X1 U625 ( .A(KEYINPUT34), .ZN(n533) );
  NOR2_X1 U626 ( .A1(n544), .A2(n542), .ZN(n591) );
  XNOR2_X1 U627 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n534) );
  OR2_X1 U628 ( .A1(n536), .A2(KEYINPUT44), .ZN(n535) );
  INV_X1 U629 ( .A(KEYINPUT88), .ZN(n536) );
  NAND2_X1 U630 ( .A1(n673), .A2(n615), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n540), .A2(n539), .ZN(n720) );
  INV_X1 U632 ( .A(n544), .ZN(n541) );
  NAND2_X1 U633 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U634 ( .A(KEYINPUT107), .B(n543), .ZN(n596) );
  INV_X1 U635 ( .A(n596), .ZN(n733) );
  NAND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n737) );
  NAND2_X1 U637 ( .A1(n733), .A2(n737), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n554), .A2(n385), .ZN(n548) );
  XOR2_X1 U639 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n549) );
  XNOR2_X1 U640 ( .A(n550), .B(n549), .ZN(n736) );
  INV_X1 U641 ( .A(n682), .ZN(n680) );
  NAND2_X1 U642 ( .A1(n676), .A2(n680), .ZN(n552) );
  INV_X1 U643 ( .A(n551), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n552), .A2(n583), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n554), .A2(n553), .ZN(n722) );
  NAND2_X1 U646 ( .A1(n736), .A2(n722), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U648 ( .A1(KEYINPUT44), .A2(n715), .ZN(n560) );
  INV_X1 U649 ( .A(KEYINPUT64), .ZN(n564) );
  NOR2_X2 U650 ( .A1(n661), .A2(n629), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT82), .ZN(n628) );
  NOR2_X1 U652 ( .A1(G900), .A2(n567), .ZN(n568) );
  NOR2_X1 U653 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U654 ( .A(KEYINPUT78), .B(n570), .ZN(n589) );
  OR2_X1 U655 ( .A1(n673), .A2(n589), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n571), .A2(n439), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n578), .A2(n385), .ZN(n573) );
  XNOR2_X1 U658 ( .A(KEYINPUT112), .B(KEYINPUT28), .ZN(n572) );
  XNOR2_X1 U659 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X1 U660 ( .A1(n574), .A2(n583), .ZN(n603) );
  NAND2_X1 U661 ( .A1(n603), .A2(n424), .ZN(n730) );
  INV_X1 U662 ( .A(n576), .ZN(n692) );
  NOR2_X1 U663 ( .A1(n730), .A2(n692), .ZN(n577) );
  XOR2_X1 U664 ( .A(KEYINPUT47), .B(n577), .Z(n581) );
  NAND2_X1 U665 ( .A1(n596), .A2(n578), .ZN(n612) );
  NOR2_X1 U666 ( .A1(n362), .A2(n615), .ZN(n579) );
  XNOR2_X1 U667 ( .A(n579), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n581), .A2(n739), .ZN(n593) );
  BUF_X2 U669 ( .A(n582), .Z(n621) );
  NOR2_X1 U670 ( .A1(n584), .A2(n583), .ZN(n588) );
  INV_X1 U671 ( .A(n613), .ZN(n687) );
  NOR2_X1 U672 ( .A1(n680), .A2(n687), .ZN(n586) );
  XNOR2_X1 U673 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n585) );
  XNOR2_X1 U674 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U675 ( .A1(n621), .A2(n594), .ZN(n590) );
  XNOR2_X1 U676 ( .A(KEYINPUT111), .B(n590), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n729) );
  NAND2_X1 U678 ( .A1(n593), .A2(n729), .ZN(n610) );
  XOR2_X1 U679 ( .A(KEYINPUT72), .B(KEYINPUT39), .Z(n595) );
  AND2_X1 U680 ( .A1(n623), .A2(n596), .ZN(n597) );
  XNOR2_X1 U681 ( .A(n597), .B(KEYINPUT40), .ZN(n780) );
  INV_X1 U682 ( .A(n780), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n605) );
  XNOR2_X1 U684 ( .A(n599), .B(KEYINPUT113), .ZN(n691) );
  NOR2_X1 U685 ( .A1(n600), .A2(n691), .ZN(n602) );
  INV_X1 U686 ( .A(KEYINPUT41), .ZN(n601) );
  XNOR2_X1 U687 ( .A(n602), .B(n601), .ZN(n704) );
  NAND2_X1 U688 ( .A1(n704), .A2(n603), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n605), .B(n604), .ZN(n778) );
  INV_X1 U690 ( .A(n778), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT48), .ZN(n627) );
  INV_X1 U693 ( .A(n612), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT43), .B(n619), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT109), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n742) );
  INV_X1 U700 ( .A(n737), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n741) );
  INV_X1 U702 ( .A(n741), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n742), .A2(n625), .ZN(n626) );
  AND2_X2 U704 ( .A1(n627), .A2(n626), .ZN(n770) );
  NAND2_X1 U705 ( .A1(n628), .A2(n770), .ZN(n632) );
  INV_X1 U706 ( .A(n629), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  INV_X1 U708 ( .A(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U709 ( .A1(n749), .A2(G472), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U711 ( .A(G952), .ZN(n638) );
  NOR2_X2 U712 ( .A1(n639), .A2(n753), .ZN(n641) );
  INV_X1 U713 ( .A(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n749), .A2(G210), .ZN(n646) );
  XOR2_X1 U716 ( .A(KEYINPUT79), .B(KEYINPUT54), .Z(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X2 U720 ( .A1(n647), .A2(n753), .ZN(n649) );
  XOR2_X1 U721 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(G51) );
  NAND2_X1 U723 ( .A1(n749), .A2(G475), .ZN(n655) );
  XOR2_X1 U724 ( .A(KEYINPUT91), .B(KEYINPUT65), .Z(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n650) );
  XOR2_X1 U726 ( .A(n651), .B(n650), .Z(n652) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U728 ( .A1(n656), .A2(n753), .ZN(n659) );
  XNOR2_X1 U729 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT66), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(G60) );
  INV_X1 U732 ( .A(KEYINPUT81), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n664), .A2(KEYINPUT81), .ZN(n665) );
  NOR2_X1 U735 ( .A1(n770), .A2(n665), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n430), .A2(n666), .ZN(n667) );
  INV_X1 U737 ( .A(KEYINPUT83), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n672), .B(n671), .ZN(n710) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n675), .Z(n679) );
  XNOR2_X1 U741 ( .A(n677), .B(KEYINPUT50), .ZN(n678) );
  OR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n547), .A2(n385), .ZN(n683) );
  NAND2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(n685), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n686), .A2(n704), .ZN(n700) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U749 ( .A1(n690), .A2(n689), .ZN(n695) );
  NOR2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U751 ( .A(KEYINPUT117), .B(n693), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT118), .ZN(n698) );
  INV_X1 U754 ( .A(n705), .ZN(n697) );
  NAND2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U757 ( .A(n701), .B(KEYINPUT52), .Z(n703) );
  NOR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n708) );
  INV_X1 U759 ( .A(n704), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n711), .B(KEYINPUT119), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n712), .A2(n771), .ZN(n714) );
  INV_X1 U765 ( .A(KEYINPUT53), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(G75) );
  XOR2_X1 U767 ( .A(n715), .B(G122), .Z(G24) );
  NAND2_X1 U768 ( .A1(n349), .A2(G217), .ZN(n718) );
  XOR2_X1 U769 ( .A(KEYINPUT123), .B(n716), .Z(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n719), .A2(n753), .ZN(G66) );
  XNOR2_X1 U772 ( .A(G101), .B(n720), .ZN(G3) );
  NOR2_X1 U773 ( .A1(n733), .A2(n722), .ZN(n721) );
  XOR2_X1 U774 ( .A(G104), .B(n721), .Z(G6) );
  NOR2_X1 U775 ( .A1(n737), .A2(n722), .ZN(n724) );
  XNOR2_X1 U776 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U778 ( .A(G107), .B(n725), .ZN(G9) );
  XNOR2_X1 U779 ( .A(G110), .B(n726), .ZN(G12) );
  NOR2_X1 U780 ( .A1(n737), .A2(n730), .ZN(n728) );
  XNOR2_X1 U781 ( .A(G128), .B(KEYINPUT29), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(G30) );
  XNOR2_X1 U783 ( .A(G143), .B(n729), .ZN(G45) );
  NOR2_X1 U784 ( .A1(n733), .A2(n730), .ZN(n732) );
  XNOR2_X1 U785 ( .A(G146), .B(KEYINPUT115), .ZN(n731) );
  XNOR2_X1 U786 ( .A(n732), .B(n731), .ZN(G48) );
  NOR2_X1 U787 ( .A1(n733), .A2(n736), .ZN(n734) );
  XOR2_X1 U788 ( .A(KEYINPUT116), .B(n734), .Z(n735) );
  XNOR2_X1 U789 ( .A(G113), .B(n735), .ZN(G15) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U791 ( .A(G116), .B(n738), .Z(G18) );
  XNOR2_X1 U792 ( .A(n739), .B(G125), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n740), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U794 ( .A(G134), .B(n741), .ZN(G36) );
  XOR2_X1 U795 ( .A(G140), .B(n742), .Z(G42) );
  NAND2_X1 U796 ( .A1(n349), .A2(G469), .ZN(n747) );
  XNOR2_X1 U797 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n743) );
  XOR2_X1 U798 ( .A(n743), .B(KEYINPUT57), .Z(n744) );
  XNOR2_X1 U799 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U801 ( .A1(n753), .A2(n748), .ZN(G54) );
  NAND2_X1 U802 ( .A1(n749), .A2(G478), .ZN(n750) );
  XOR2_X1 U803 ( .A(n751), .B(n750), .Z(n752) );
  NOR2_X1 U804 ( .A1(n753), .A2(n752), .ZN(G63) );
  NOR2_X1 U805 ( .A1(n754), .A2(G953), .ZN(n760) );
  NAND2_X1 U806 ( .A1(G224), .A2(G953), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n755), .B(KEYINPUT124), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n757), .A2(n761), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n758), .B(KEYINPUT125), .ZN(n759) );
  NOR2_X1 U811 ( .A1(n760), .A2(n759), .ZN(n767) );
  NOR2_X1 U812 ( .A1(n761), .A2(n771), .ZN(n765) );
  XOR2_X1 U813 ( .A(G101), .B(G110), .Z(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U815 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U816 ( .A(n767), .B(n766), .Z(G69) );
  XOR2_X1 U817 ( .A(n768), .B(n769), .Z(n773) );
  XNOR2_X1 U818 ( .A(n770), .B(n773), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(n771), .ZN(n777) );
  XOR2_X1 U820 ( .A(G227), .B(n773), .Z(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U824 ( .A(n778), .B(G137), .Z(G39) );
  XOR2_X1 U825 ( .A(G131), .B(KEYINPUT126), .Z(n779) );
  XNOR2_X1 U826 ( .A(n780), .B(n779), .ZN(G33) );
  XNOR2_X1 U827 ( .A(n781), .B(G119), .ZN(G21) );
endmodule

