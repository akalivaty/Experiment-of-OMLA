//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G244), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n214), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n250), .A2(new_n252), .B1(G50), .B2(new_n249), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n215), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n201), .A2(new_n215), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n246), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n255), .A2(KEYINPUT74), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT74), .B1(new_n255), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT9), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n255), .A2(new_n263), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  AND4_X1   g0083(.A1(new_n277), .A2(new_n279), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G223), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(G1698), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n202), .B2(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  INV_X1    g0093(.A(new_n214), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n291), .A3(G274), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT66), .B(G226), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n297), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  MUX2_X1   g0110(.A(new_n274), .B(new_n275), .S(new_n310), .Z(new_n311));
  NAND2_X1  g0111(.A1(new_n273), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n273), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n277), .A2(new_n279), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G107), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n277), .A2(new_n279), .A3(new_n281), .A4(new_n283), .ZN(new_n319));
  INV_X1    g0119(.A(G238), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n318), .B1(new_n319), .B2(new_n233), .C1(new_n320), .C2(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n296), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n307), .A2(new_n218), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n301), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n256), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT15), .B(G87), .Z(new_n329));
  INV_X1    g0129(.A(new_n257), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n246), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  INV_X1    g0134(.A(new_n249), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n202), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n246), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G77), .A3(new_n251), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n334), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n247), .B1(new_n328), .B2(new_n331), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n336), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT72), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n326), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n324), .A2(G179), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n326), .A2(new_n343), .A3(KEYINPUT73), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(G200), .B2(new_n324), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n274), .B2(new_n324), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n310), .A2(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n310), .A2(new_n325), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n268), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT71), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n316), .A2(new_n349), .A3(new_n351), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n330), .A2(G77), .B1(G20), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G50), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n260), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT11), .A3(new_n246), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n337), .A2(G68), .A3(new_n251), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT77), .B1(new_n335), .B2(new_n357), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n360), .A2(new_n246), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n363), .B(new_n365), .C1(KEYINPUT11), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n281), .A2(new_n283), .A3(G226), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G232), .A2(G1698), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n317), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n296), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT67), .B1(new_n291), .B2(new_n302), .ZN(new_n376));
  OAI21_X1  g0176(.A(G238), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n373), .A2(new_n374), .A3(new_n301), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n291), .A2(G274), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n307), .A2(G238), .B1(new_n381), .B2(new_n300), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n374), .A4(new_n373), .ZN(new_n384));
  INV_X1    g0184(.A(new_n373), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n377), .A2(new_n301), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT13), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n379), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G169), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(G179), .A3(new_n378), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n388), .B2(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n367), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n367), .B1(new_n388), .B2(G200), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(G190), .A3(new_n378), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n387), .A2(KEYINPUT76), .A3(G190), .A4(new_n378), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n327), .A2(new_n251), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n250), .B1(new_n249), .B2(new_n327), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n286), .B2(G20), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(G20), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n317), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n357), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  AND2_X1   g0212(.A1(G58), .A2(G68), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G58), .A2(G68), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(G20), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n259), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(G58), .B(G68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n418), .B2(G20), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT79), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(G20), .B1(new_n413), .B2(new_n414), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT79), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n416), .A4(new_n415), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n411), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n247), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n276), .A2(KEYINPUT80), .A3(G33), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n409), .B(new_n428), .C1(new_n317), .C2(KEYINPUT80), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n357), .B1(new_n429), .B2(new_n408), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n416), .A3(new_n415), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n406), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n291), .A2(G232), .A3(new_n302), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT83), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n301), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n301), .B2(new_n434), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G87), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n319), .A2(new_n287), .B1(new_n278), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT82), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n286), .A2(new_n441), .A3(G226), .A4(G1698), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n277), .A2(new_n279), .A3(G226), .A4(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n291), .B(KEYINPUT69), .ZN(new_n446));
  OAI211_X1 g0246(.A(G179), .B(new_n438), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n278), .A2(new_n439), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n284), .B2(G223), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n442), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n301), .A2(new_n434), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n301), .A2(new_n434), .A3(new_n435), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G169), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT18), .B1(new_n433), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n274), .B(new_n438), .C1(new_n445), .C2(new_n446), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n275), .B1(new_n451), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n420), .A2(new_n424), .ZN(new_n462));
  INV_X1    g0262(.A(new_n411), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(KEYINPUT16), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n246), .A3(new_n432), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n404), .B(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n466), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n447), .A2(new_n456), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n461), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n458), .A2(new_n469), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n356), .A2(new_n402), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT68), .B(G1698), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n286), .A2(new_n477), .A3(KEYINPUT4), .A4(G244), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT4), .B1(new_n284), .B2(G244), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n296), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n299), .A2(G1), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n380), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n291), .ZN(new_n490));
  INV_X1    g0290(.A(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n487), .A2(KEYINPUT85), .A3(G257), .A4(new_n291), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G179), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n483), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(new_n494), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n325), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n499), .A2(new_n204), .A3(G107), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n502), .A2(new_n215), .B1(new_n202), .B2(new_n260), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n205), .B1(new_n429), .B2(new_n408), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(KEYINPUT84), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n429), .A2(new_n408), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G107), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n247), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n249), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n248), .A2(G33), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n214), .A2(new_n249), .A3(new_n245), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(G97), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n496), .B(new_n498), .C1(new_n510), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n506), .A2(KEYINPUT84), .A3(G107), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n499), .ZN(new_n518));
  INV_X1    g0318(.A(new_n500), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n246), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n483), .A2(new_n494), .A3(new_n274), .ZN(new_n525));
  AOI21_X1  g0325(.A(G200), .B1(new_n483), .B2(new_n494), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n514), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n329), .A2(new_n249), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n215), .B1(new_n371), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G87), .B2(new_n206), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n277), .A2(new_n279), .A3(new_n215), .A4(G68), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n257), .B2(new_n204), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n528), .B1(new_n534), .B2(new_n246), .ZN(new_n535));
  INV_X1    g0335(.A(new_n329), .ZN(new_n536));
  INV_X1    g0336(.A(new_n513), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n484), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n291), .ZN(new_n541));
  INV_X1    g0341(.A(new_n484), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n380), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n277), .A2(new_n279), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n319), .C2(new_n320), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n296), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n325), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n296), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n381), .A2(new_n484), .B1(new_n291), .B2(new_n540), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n549), .A2(G179), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n538), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n535), .B1(new_n439), .B2(new_n537), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n275), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT86), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI221_X4 g0355(.A(new_n528), .B1(new_n513), .B2(G87), .C1(new_n534), .C2(new_n246), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n275), .C2(new_n547), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n547), .A2(G190), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND4_X1   g0360(.A1(new_n516), .A2(new_n527), .A3(new_n552), .A4(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n277), .A2(new_n279), .A3(new_n215), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n286), .A2(new_n564), .A3(new_n215), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n545), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n215), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n566), .A2(new_n573), .A3(new_n571), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n247), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT89), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT25), .ZN(new_n579));
  AOI21_X1  g0379(.A(G107), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n335), .A2(new_n580), .B1(KEYINPUT89), .B2(KEYINPUT25), .ZN(new_n581));
  NOR4_X1   g0381(.A1(new_n249), .A2(new_n578), .A3(new_n579), .A4(G107), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n537), .A2(new_n205), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n277), .A2(new_n279), .A3(G257), .A4(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G294), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n319), .C2(new_n539), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n296), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n380), .A2(new_n487), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n487), .A2(new_n291), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G264), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(new_n274), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT90), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n275), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n587), .A2(new_n296), .B1(new_n590), .B2(G264), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT90), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(new_n274), .A4(new_n589), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n584), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n495), .A3(new_n589), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n594), .A2(new_n325), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n577), .C2(new_n583), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n286), .A2(new_n477), .A3(G257), .ZN(new_n605));
  XOR2_X1   g0405(.A(KEYINPUT87), .B(G303), .Z(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n286), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G264), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n288), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n296), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n488), .B1(new_n590), .B2(G270), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n513), .A2(G116), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n335), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n245), .A2(new_n214), .B1(G20), .B2(new_n614), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n480), .B(new_n215), .C1(G33), .C2(new_n204), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n616), .A2(KEYINPUT20), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT20), .B1(new_n616), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n613), .B(new_n615), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n612), .A2(G169), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n620), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n610), .A2(G190), .A3(new_n611), .ZN(new_n625));
  INV_X1    g0425(.A(G270), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n589), .B1(new_n626), .B2(new_n490), .ZN(new_n627));
  OAI221_X1 g0427(.A(new_n605), .B1(new_n286), .B2(new_n606), .C1(new_n608), .C2(new_n288), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n296), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n624), .B(new_n625), .C1(new_n629), .C2(new_n275), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(G179), .A3(new_n620), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n612), .A2(KEYINPUT21), .A3(G169), .A4(new_n620), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n623), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n604), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n476), .A2(new_n561), .A3(new_n634), .ZN(G372));
  OAI21_X1  g0435(.A(KEYINPUT91), .B1(new_n548), .B2(new_n551), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n547), .A2(G179), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT91), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n325), .C2(new_n547), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n538), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n553), .A2(new_n554), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n640), .A2(new_n538), .B1(new_n642), .B2(new_n559), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n631), .A2(new_n632), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n603), .A3(new_n623), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n645), .A3(new_n600), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n516), .A2(new_n527), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n560), .A2(new_n552), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n649), .A2(new_n650), .A3(new_n516), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n516), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n524), .A2(new_n514), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT92), .A3(new_n496), .A4(new_n498), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n643), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n656), .B2(new_n650), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n476), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n355), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n348), .A2(new_n347), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT73), .B1(new_n326), .B2(new_n343), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT93), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT93), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n346), .A2(new_n664), .A3(new_n347), .A4(new_n348), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n388), .A2(G169), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT14), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n391), .A3(new_n390), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n663), .A2(new_n665), .B1(new_n668), .B2(new_n367), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n401), .A2(new_n469), .A3(new_n474), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n458), .B(new_n473), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n660), .B1(new_n671), .B2(new_n316), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n659), .A2(new_n672), .ZN(G369));
  NAND2_X1  g0473(.A1(new_n644), .A2(new_n623), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n248), .A2(new_n215), .A3(G13), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT94), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G213), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n624), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n674), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n633), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n685), .A2(new_n584), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n604), .A2(new_n691), .B1(new_n603), .B2(new_n685), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n674), .A2(new_n685), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(new_n604), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n603), .B2(new_n684), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n694), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n212), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n705));
  XNOR2_X1  g0505(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n658), .A2(new_n685), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n516), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n552), .A3(new_n560), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n641), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(KEYINPUT26), .B2(new_n656), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n647), .B(KEYINPUT97), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n643), .A2(new_n600), .A3(new_n645), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n714), .A2(KEYINPUT98), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT98), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n483), .A2(new_n494), .A3(new_n547), .A4(new_n596), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n610), .A2(G179), .A3(new_n611), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n483), .A2(new_n494), .A3(new_n547), .A4(new_n596), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT30), .B1(new_n727), .B2(new_n724), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n629), .A2(G179), .A3(new_n547), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n497), .A2(new_n594), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n726), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n684), .A2(KEYINPUT31), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n731), .A2(KEYINPUT96), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT96), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n634), .A2(new_n561), .A3(new_n685), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n731), .B2(new_n685), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(G330), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n721), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT99), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n706), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n248), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n700), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n690), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G330), .B2(new_n688), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n286), .A2(new_n209), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n209), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n317), .A2(new_n209), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT100), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n299), .B2(new_n213), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n240), .A2(new_n299), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n214), .B1(G20), .B2(new_n325), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n748), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n215), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n495), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n317), .B1(new_n768), .B2(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n215), .A2(new_n275), .A3(G179), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n215), .B1(new_n767), .B2(G190), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n215), .A2(new_n495), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT101), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT101), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n773), .B(new_n779), .C1(new_n785), .C2(G326), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n274), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n780), .A2(new_n274), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G317), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n771), .A2(G20), .A3(G190), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n791), .A2(G283), .B1(new_n800), .B2(KEYINPUT103), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n786), .B(new_n801), .C1(KEYINPUT103), .C2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n790), .A2(new_n205), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G50), .B2(new_n785), .ZN(new_n804));
  INV_X1    g0604(.A(new_n768), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G159), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G68), .B2(new_n793), .ZN(new_n808));
  INV_X1    g0608(.A(G58), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n286), .B1(new_n772), .B2(new_n202), .C1(new_n809), .C2(new_n799), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n778), .A2(new_n204), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n775), .A2(new_n439), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n804), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n802), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n765), .B1(new_n815), .B2(new_n762), .ZN(new_n816));
  INV_X1    g0616(.A(new_n761), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n688), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n750), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n684), .A2(new_n343), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n663), .A2(new_n665), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n349), .A2(new_n351), .A3(new_n821), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n707), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n685), .C1(new_n648), .C2(new_n657), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n748), .B1(new_n829), .B2(new_n740), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n740), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n762), .A2(new_n759), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT104), .Z(new_n833));
  OAI21_X1  g0633(.A(new_n748), .B1(new_n833), .B2(G77), .ZN(new_n834));
  INV_X1    g0634(.A(new_n799), .ZN(new_n835));
  INV_X1    g0635(.A(new_n772), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G294), .B1(new_n836), .B2(G116), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n770), .B2(new_n768), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n811), .B(new_n838), .C1(G283), .C2(new_n793), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n317), .B1(new_n775), .B2(new_n205), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT105), .Z(new_n841));
  NAND2_X1  g0641(.A1(new_n791), .A2(G87), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n785), .A2(G303), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n791), .A2(G68), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n286), .B1(new_n846), .B2(new_n768), .C1(new_n775), .C2(new_n359), .ZN(new_n847));
  INV_X1    g0647(.A(new_n778), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(G58), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n835), .A2(G143), .B1(new_n836), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n258), .B2(new_n792), .C1(new_n784), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n845), .B(new_n849), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n852), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n834), .B1(new_n857), .B2(new_n762), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n825), .B2(new_n760), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n831), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n745), .A2(new_n248), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n395), .A2(new_n400), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n367), .B(new_n684), .C1(new_n863), .C2(new_n668), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n367), .A2(new_n684), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n394), .A2(new_n401), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n462), .A2(new_n463), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n427), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n406), .B1(new_n426), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n467), .B1(new_n870), .B2(new_n682), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n457), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n470), .A2(new_n472), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n470), .A2(new_n681), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n467), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n870), .A2(new_n682), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n475), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n349), .A2(new_n684), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n828), .A2(KEYINPUT106), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT106), .B1(new_n828), .B2(new_n884), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n867), .B1(new_n881), .B2(new_n882), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n681), .B1(new_n458), .B2(new_n473), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT107), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n467), .B1(new_n433), .B2(new_n457), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n433), .A2(new_n682), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n877), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n475), .A2(new_n892), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT107), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n878), .A2(new_n880), .A3(new_n900), .A4(KEYINPUT38), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n890), .A2(new_n898), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n882), .A2(new_n881), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n668), .A2(new_n367), .A3(new_n685), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n888), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n887), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n709), .A2(new_n719), .A3(new_n476), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n672), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n908), .B(new_n910), .Z(new_n911));
  NAND2_X1  g0711(.A1(new_n726), .A2(new_n728), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n729), .A2(new_n730), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT109), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT31), .A4(new_n684), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT109), .B1(new_n731), .B2(new_n732), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n736), .A2(new_n738), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  AND4_X1   g0718(.A1(KEYINPUT40), .A2(new_n867), .A3(new_n918), .A4(new_n825), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n890), .A2(new_n901), .A3(new_n898), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n867), .A2(new_n918), .A3(new_n825), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n903), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n476), .A2(new_n918), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(G330), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n862), .B1(new_n911), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n911), .B2(new_n930), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(G116), .A3(new_n216), .A4(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n212), .A2(new_n413), .A3(new_n202), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n357), .A2(G50), .ZN(new_n938));
  OAI211_X1 g0738(.A(G1), .B(new_n744), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n936), .A3(new_n939), .ZN(G367));
  NOR2_X1   g0740(.A1(new_n231), .A2(new_n755), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n763), .B1(new_n209), .B2(new_n536), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n748), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n791), .A2(G77), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n785), .A2(G143), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n772), .A2(new_n359), .B1(new_n768), .B2(new_n851), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n317), .B(new_n946), .C1(G150), .C2(new_n835), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n778), .A2(new_n357), .ZN(new_n948));
  INV_X1    g0748(.A(G159), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n792), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n775), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n948), .B(new_n950), .C1(G58), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n944), .A2(new_n945), .A3(new_n947), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n791), .A2(G97), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n784), .B2(new_n770), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(G116), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  INV_X1    g0757(.A(G283), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n772), .A2(new_n958), .B1(new_n768), .B2(new_n794), .ZN(new_n959));
  INV_X1    g0759(.A(new_n606), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n286), .B(new_n959), .C1(new_n960), .C2(new_n835), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n793), .A2(G294), .B1(new_n848), .B2(G107), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n957), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n953), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n943), .B1(new_n965), .B2(new_n762), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n643), .B1(new_n556), .B2(new_n685), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n640), .A2(new_n538), .A3(new_n553), .A4(new_n684), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n969), .B2(new_n817), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n654), .A2(new_n684), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n714), .A2(new_n972), .B1(new_n710), .B2(new_n684), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n696), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT42), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n973), .B(KEYINPUT110), .Z(new_n977));
  INV_X1    g0777(.A(new_n603), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n710), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n971), .B(new_n976), .C1(new_n979), .C2(new_n684), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT111), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n969), .B(KEYINPUT43), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n979), .A2(new_n684), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n975), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n694), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n982), .A2(new_n694), .A3(new_n977), .A4(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n973), .A2(new_n697), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT112), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n973), .A2(new_n697), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT45), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(new_n694), .ZN(new_n999));
  INV_X1    g0799(.A(new_n695), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n696), .B1(new_n692), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(new_n689), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n742), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n700), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n747), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n970), .B1(new_n990), .B2(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(new_n1002), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n692), .A2(new_n817), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n751), .A2(new_n702), .B1(G107), .B2(new_n209), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n236), .A2(new_n299), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n702), .B(new_n299), .C1(new_n357), .C2(new_n202), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n256), .B2(G50), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n327), .A2(KEYINPUT50), .A3(new_n359), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n755), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1010), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n748), .B1(new_n1018), .B2(new_n764), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n775), .A2(new_n202), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n536), .A2(new_n778), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n327), .C2(new_n793), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n772), .A2(new_n357), .B1(new_n768), .B2(new_n258), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n317), .B(new_n1023), .C1(G50), .C2(new_n835), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n785), .A2(G159), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n954), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n286), .B1(new_n805), .B2(G326), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n775), .A2(new_n777), .B1(new_n958), .B2(new_n778), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n836), .A2(new_n960), .B1(new_n835), .B2(G317), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n770), .B2(new_n792), .C1(new_n784), .C2(new_n798), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1027), .B1(new_n614), .B2(new_n790), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1019), .B1(new_n1037), .B2(new_n762), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1008), .A2(new_n747), .B1(new_n1009), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n742), .A2(new_n1008), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n700), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n742), .A2(new_n1008), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  XNOR2_X1  g0843(.A(new_n998), .B(new_n693), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n747), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n763), .B1(new_n204), .B2(new_n209), .C1(new_n755), .C2(new_n243), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n748), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n784), .A2(new_n258), .B1(new_n949), .B2(new_n799), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n775), .A2(new_n357), .B1(new_n202), .B2(new_n778), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n317), .B1(new_n805), .B2(G143), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n256), .B2(new_n772), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G50), .C2(new_n793), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n842), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n784), .A2(new_n794), .B1(new_n770), .B2(new_n799), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n951), .A2(G283), .B1(new_n848), .B2(G116), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n606), .B2(new_n792), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n317), .B1(new_n768), .B2(new_n798), .C1(new_n777), .C2(new_n772), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n803), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1047), .B1(new_n1061), .B2(new_n762), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n977), .B2(new_n817), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n700), .B1(new_n1040), .B2(new_n999), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1044), .B1(new_n742), .B2(new_n1008), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1045), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  NAND4_X1  g0866(.A1(new_n867), .A2(new_n918), .A3(G330), .A4(new_n825), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n867), .B1(new_n885), .B2(new_n886), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n904), .B1(new_n1069), .B2(new_n905), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n920), .A2(new_n905), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n718), .A2(new_n685), .A3(new_n825), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n884), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1073), .B2(new_n867), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT113), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n927), .A2(G330), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n672), .A3(new_n909), .ZN(new_n1078));
  OAI211_X1 g0878(.A(G330), .B(new_n825), .C1(new_n735), .C2(new_n739), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n867), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1067), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n885), .B2(new_n886), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT114), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(KEYINPUT114), .C1(new_n886), .C2(new_n885), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n918), .A2(G330), .A3(new_n825), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1080), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1088), .A2(new_n1072), .A3(new_n884), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1078), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1088), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT113), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n1068), .C1(new_n1070), .C2(new_n1074), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1076), .A2(new_n1092), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1092), .B(KEYINPUT115), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1076), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n700), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n904), .A2(new_n760), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n748), .B1(new_n833), .B2(new_n327), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n799), .A2(new_n614), .B1(new_n772), .B2(new_n204), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n286), .B(new_n1103), .C1(G294), .C2(new_n805), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n785), .A2(G283), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n778), .A2(new_n202), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1106), .B(new_n812), .C1(G107), .C2(new_n793), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n845), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n775), .A2(new_n258), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n317), .B1(new_n836), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n835), .A2(G132), .B1(new_n805), .B2(G125), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n793), .A2(G137), .B1(new_n848), .B2(G159), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n790), .A2(new_n359), .B1(new_n784), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1102), .B1(new_n1118), .B2(new_n762), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1099), .A2(new_n747), .B1(new_n1101), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1100), .A2(new_n1120), .ZN(G378));
  INV_X1    g0921(.A(new_n1078), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n921), .A2(new_n925), .A3(G330), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n682), .B1(new_n270), .B2(new_n264), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n316), .B2(new_n354), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n354), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1131), .B(new_n1128), .C1(new_n313), .C2(new_n315), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n315), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n314), .B1(new_n273), .B2(new_n311), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n354), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1128), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n316), .A2(new_n354), .A3(new_n1129), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1126), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1124), .A2(new_n1125), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1125), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n921), .A3(new_n925), .A4(G330), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n908), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT117), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n887), .A2(new_n1145), .A3(new_n907), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1143), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT116), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1124), .A2(new_n1140), .A3(new_n1125), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n887), .A2(new_n1145), .A3(new_n907), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT117), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1147), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1123), .A2(new_n1157), .A3(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1097), .A2(new_n1122), .B1(new_n1147), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n700), .C1(KEYINPUT57), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1140), .A2(new_n759), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n832), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n748), .B1(G50), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n359), .B1(G33), .B2(G41), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n317), .B2(new_n298), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n791), .A2(G58), .B1(new_n785), .B2(G116), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G41), .B(new_n286), .C1(new_n805), .C2(G283), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n835), .A2(G107), .B1(new_n836), .B2(new_n329), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n948), .B(new_n1020), .C1(G97), .C2(new_n793), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n799), .A2(new_n1116), .B1(new_n772), .B2(new_n851), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G132), .B2(new_n793), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n951), .A2(new_n1111), .B1(new_n848), .B2(G150), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1176), .C1(new_n1177), .C2(new_n784), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n949), .C2(new_n790), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1179), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1164), .B1(new_n1183), .B2(new_n762), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1162), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1147), .A2(new_n1159), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n747), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1161), .A2(new_n1188), .ZN(G375));
  NAND2_X1  g0989(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1080), .A2(new_n759), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n748), .B1(new_n833), .B2(G68), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n286), .B1(new_n768), .B2(new_n1116), .C1(new_n258), .C2(new_n772), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n775), .A2(new_n949), .B1(new_n359), .B2(new_n778), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n791), .C2(G58), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT119), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n793), .A2(new_n1111), .B1(new_n835), .B2(G137), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n784), .A2(new_n846), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(KEYINPUT118), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(KEYINPUT118), .B2(new_n1198), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n792), .A2(new_n614), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1202), .B(new_n1021), .C1(G97), .C2(new_n951), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n799), .A2(new_n958), .B1(new_n772), .B2(new_n205), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n286), .B(new_n1204), .C1(G303), .C2(new_n805), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n785), .A2(G294), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n944), .A2(new_n1203), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1192), .B1(new_n1208), .B2(new_n762), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1190), .A2(new_n747), .B1(new_n1191), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1087), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1005), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1098), .B2(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G390), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n860), .ZN(new_n1215));
  OR2_X1    g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(new_n1216), .A3(G387), .A4(G381), .ZN(new_n1217));
  INV_X1    g1017(.A(G378), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1161), .A4(new_n1188), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n683), .A2(G213), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G407), .B(G213), .C1(G375), .C2(new_n1222), .ZN(G409));
  INV_X1    g1023(.A(KEYINPUT122), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1160), .A2(new_n1005), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n746), .B1(new_n1157), .B2(KEYINPUT120), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1148), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1154), .A2(KEYINPUT117), .A3(new_n1155), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1154), .A2(new_n1145), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1227), .A2(new_n1228), .B1(new_n1229), .B2(new_n908), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT120), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1186), .B1(new_n1226), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1225), .B1(new_n1233), .B2(KEYINPUT121), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n747), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1185), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT121), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G378), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1161), .A2(G378), .A3(new_n1188), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1224), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1190), .A2(new_n1122), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT60), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(new_n1211), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1211), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n700), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1210), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n860), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(G384), .A3(new_n1210), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(KEYINPUT121), .B(new_n1185), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1160), .A2(new_n1005), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1226), .A2(new_n1232), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT121), .B1(new_n1256), .B2(new_n1185), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1218), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1161), .A2(G378), .A3(new_n1188), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(KEYINPUT122), .A3(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1242), .A2(new_n1220), .A3(new_n1252), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n990), .A2(new_n1006), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n970), .A3(G390), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1214), .A2(G387), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n819), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1221), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1251), .A2(new_n1262), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1276), .B2(KEYINPUT123), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1242), .A2(new_n1220), .A3(new_n1260), .ZN(new_n1278));
  INV_X1    g1078(.A(G2897), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1251), .A2(new_n1279), .A3(new_n1220), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1249), .A2(new_n1250), .B1(G2897), .B2(new_n1221), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1274), .A2(new_n1285), .A3(new_n1275), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1263), .A2(new_n1277), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1271), .B1(new_n1282), .B2(new_n1274), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1261), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1274), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(new_n1259), .A2(KEYINPUT124), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1218), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1295), .B(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1251), .B2(KEYINPUT125), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1298), .B2(new_n1251), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1293), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1293), .A2(new_n1303), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1299), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1302), .A2(new_n1304), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1303), .B(new_n1293), .C1(new_n1309), .C2(new_n1301), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(G402));
endmodule


