//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  AOI21_X1  g005(.A(G107), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(G101), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NOR3_X1   g009(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n192), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(new_n191), .A3(G107), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT64), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G146), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G143), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT64), .B(G143), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(new_n209), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT80), .B(new_n195), .C1(new_n199), .C2(new_n202), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n205), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT10), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n210), .ZN(new_n224));
  AOI21_X1  g038(.A(G146), .B1(new_n206), .B2(new_n207), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(G128), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n222), .B1(new_n228), .B2(new_n203), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n208), .A2(new_n210), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT64), .A2(G143), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT64), .A2(G143), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n211), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n213), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT77), .B(G104), .ZN(new_n237));
  AOI21_X1  g051(.A(G101), .B1(new_n237), .B2(G107), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(new_n197), .C1(new_n198), .C2(new_n192), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n236), .A2(new_n239), .A3(KEYINPUT79), .A4(new_n195), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n229), .A2(new_n230), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n221), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT11), .A3(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n245), .A2(new_n247), .A3(new_n251), .A4(new_n248), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n200), .B(new_n197), .C1(new_n192), .C2(new_n198), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G101), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n225), .B2(new_n214), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n208), .A2(new_n210), .A3(new_n257), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n239), .A3(KEYINPUT4), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n190), .A2(G104), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n193), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n196), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n255), .B1(new_n270), .B2(new_n238), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT78), .B1(new_n271), .B2(new_n263), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n262), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n242), .A2(new_n253), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n218), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n229), .A2(new_n240), .B1(new_n275), .B2(new_n203), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT12), .B1(new_n276), .B2(new_n253), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n250), .A2(new_n252), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n229), .A2(new_n240), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n218), .B1(new_n239), .B2(new_n195), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G110), .B(G140), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n284), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n242), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n279), .ZN(new_n290));
  INV_X1    g104(.A(new_n287), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n274), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n187), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT81), .B(G469), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n290), .B2(new_n274), .ZN(new_n297));
  AND4_X1   g111(.A1(new_n274), .A2(new_n277), .A3(new_n282), .A4(new_n291), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n294), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT82), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n242), .A2(new_n253), .A3(new_n273), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n253), .B1(new_n242), .B2(new_n273), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n287), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n274), .A2(new_n277), .A3(new_n282), .A4(new_n291), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n296), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n295), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT76), .ZN(new_n310));
  OAI21_X1  g124(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n313));
  INV_X1    g127(.A(G237), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n314), .A2(new_n285), .A3(G214), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G143), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n215), .B2(new_n315), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(G131), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G146), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n320), .A2(new_n322), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT19), .Z(new_n327));
  OAI211_X1 g141(.A(new_n318), .B(new_n325), .C1(G146), .C2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(KEYINPUT18), .A3(G131), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n326), .B(new_n209), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT18), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n251), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n329), .B(new_n330), .C1(new_n317), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G113), .B(G122), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(new_n188), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n317), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n323), .A2(G146), .A3(new_n324), .ZN(new_n340));
  AOI21_X1  g154(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n342), .A3(KEYINPUT90), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n318), .B2(KEYINPUT17), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT90), .B1(new_n339), .B2(new_n342), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n336), .B(new_n333), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G475), .A2(G902), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n313), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n313), .A3(new_n348), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n333), .B1(new_n344), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n337), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n346), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n294), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT91), .B(G475), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n350), .A2(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(G234), .A2(G237), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(G952), .A3(new_n285), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(G902), .A3(G953), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT21), .B(G898), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G478), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT15), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n310), .A2(new_n367), .A3(G953), .ZN(new_n368));
  AND2_X1   g182(.A1(KEYINPUT68), .A2(G116), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT68), .A2(G116), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G122), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G107), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n372), .B(new_n193), .C1(new_n373), .C2(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n206), .A2(G128), .A3(new_n207), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n244), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G143), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n378), .B1(G128), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(new_n380), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n378), .B(new_n244), .C1(G128), .C2(new_n382), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n385), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n390));
  OAI21_X1  g204(.A(G107), .B1(new_n372), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n388), .B(new_n376), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n368), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n392), .A3(new_n368), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n366), .B1(new_n396), .B2(new_n294), .ZN(new_n397));
  INV_X1    g211(.A(new_n395), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n294), .B(new_n366), .C1(new_n398), .C2(new_n393), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n357), .A2(new_n363), .A3(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n308), .A2(new_n312), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n404));
  INV_X1    g218(.A(G119), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(G128), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(G128), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G119), .B(G128), .ZN(new_n410));
  INV_X1    g224(.A(G110), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT24), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT24), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G110), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n409), .A2(G110), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n340), .B2(new_n341), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n409), .A2(G110), .B1(new_n410), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n326), .A2(new_n209), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n325), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G137), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n294), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT71), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT71), .B1(new_n417), .B2(new_n420), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT72), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n417), .A2(new_n420), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT71), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(KEYINPUT72), .A3(new_n435), .A4(new_n430), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT25), .B(new_n426), .C1(new_n431), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n435), .A3(new_n430), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n425), .B1(new_n443), .B2(new_n436), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT74), .B(KEYINPUT25), .Z(new_n446));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI211_X1 g262(.A(KEYINPUT73), .B(new_n425), .C1(new_n443), .C2(new_n436), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n440), .B(new_n445), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n367), .B1(G234), .B2(new_n294), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n431), .A2(new_n437), .ZN(new_n453));
  INV_X1    g267(.A(new_n424), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n451), .A2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT2), .B(G113), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n405), .A2(G116), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n371), .B2(G119), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(new_n463), .B2(KEYINPUT67), .ZN(new_n464));
  OR2_X1    g278(.A1(KEYINPUT68), .A2(G116), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT68), .A2(G116), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(G119), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n459), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n244), .A2(G137), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n246), .A2(G134), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(G131), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G134), .B(G137), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT66), .B1(new_n476), .B2(new_n251), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n218), .A2(new_n252), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n279), .A2(new_n260), .A3(new_n261), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(KEYINPUT30), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n252), .A3(new_n475), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n234), .B1(G143), .B2(new_n209), .ZN(new_n482));
  INV_X1    g296(.A(new_n217), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n484), .B2(new_n213), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n260), .A2(new_n261), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n253), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n279), .A2(KEYINPUT65), .A3(new_n260), .A4(new_n261), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n471), .B(new_n480), .C1(new_n490), .C2(KEYINPUT30), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n478), .A2(new_n479), .ZN(new_n492));
  INV_X1    g306(.A(new_n471), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n314), .A2(new_n285), .A3(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT31), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n492), .B2(new_n493), .ZN(new_n502));
  AND4_X1   g316(.A1(new_n501), .A2(new_n493), .A3(new_n478), .A4(new_n479), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n502), .A2(new_n503), .B1(new_n493), .B2(new_n490), .ZN(new_n504));
  INV_X1    g318(.A(new_n498), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n507));
  NAND4_X1  g321(.A1(new_n491), .A2(new_n494), .A3(new_n498), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n500), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G472), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n294), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT32), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n513), .A3(new_n510), .A4(new_n294), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n502), .A2(new_n503), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n492), .A2(new_n493), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT29), .A3(new_n498), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n491), .A2(new_n494), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n505), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(KEYINPUT70), .A3(new_n505), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n504), .B2(new_n505), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n294), .B(new_n519), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G472), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n458), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G214), .B1(G237), .B2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n471), .A2(new_n256), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n264), .A2(new_n265), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n271), .A2(KEYINPUT78), .A3(new_n263), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n467), .A2(KEYINPUT5), .A3(new_n461), .ZN(new_n536));
  OAI21_X1  g350(.A(G113), .B1(new_n461), .B2(KEYINPUT5), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n536), .A2(new_n538), .B1(new_n463), .B2(new_n460), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n205), .A2(new_n219), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G110), .B(G122), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n535), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n203), .A2(new_n539), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n542), .B(KEYINPUT8), .Z(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n537), .B1(new_n536), .B2(KEYINPUT85), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n463), .A2(new_n550), .A3(KEYINPUT5), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n463), .A2(new_n460), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n203), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT86), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n218), .A2(new_n321), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n260), .A2(G125), .A3(new_n261), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n285), .A2(G224), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(KEYINPUT87), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n556), .A2(new_n557), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n546), .B1(new_n203), .B2(new_n539), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n549), .A2(new_n551), .B1(new_n460), .B2(new_n463), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n567), .C1(new_n203), .C2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n555), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n294), .B1(new_n544), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT88), .B(new_n294), .C1(new_n544), .C2(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n532), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n266), .B2(new_n272), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT83), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n540), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT83), .B1(new_n535), .B2(new_n541), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n543), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT6), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n535), .A2(new_n541), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n542), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n559), .B(KEYINPUT84), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n558), .B(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n543), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n575), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n575), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n531), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n575), .A2(new_n589), .ZN(new_n596));
  INV_X1    g410(.A(new_n590), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n575), .A2(new_n589), .A3(new_n590), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(KEYINPUT89), .A3(new_n531), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n403), .A2(new_n530), .A3(new_n595), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n509), .A2(new_n294), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n452), .A2(new_n605), .A3(new_n511), .A4(new_n457), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n308), .A2(new_n606), .A3(new_n312), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n531), .B(new_n363), .C1(new_n591), .C2(new_n592), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n294), .B1(new_n398), .B2(new_n393), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n364), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n396), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n394), .A2(new_n611), .A3(new_n612), .A4(new_n395), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n294), .A2(G478), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n610), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n355), .A2(new_n356), .ZN(new_n621));
  INV_X1    g435(.A(new_n351), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n349), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n608), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n607), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(new_n401), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n357), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n608), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n607), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n605), .A2(new_n511), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT94), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT93), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n430), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n429), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n456), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n637), .B1(new_n452), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n641), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT93), .B(new_n643), .C1(new_n450), .C2(new_n451), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n636), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n451), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n443), .A2(new_n436), .ZN(new_n647));
  AND4_X1   g461(.A1(KEYINPUT75), .A2(new_n647), .A3(KEYINPUT25), .A4(new_n426), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT75), .B1(new_n444), .B2(KEYINPUT25), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT73), .B1(new_n453), .B2(new_n425), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n444), .A2(new_n447), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n652), .A3(new_n446), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n646), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT93), .B1(new_n654), .B2(new_n643), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n452), .A2(new_n637), .A3(new_n641), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(KEYINPUT94), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n635), .B1(new_n645), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n595), .A2(new_n601), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n403), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n645), .A2(new_n657), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n593), .A2(new_n308), .A3(new_n312), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n512), .A2(new_n514), .B1(new_n528), .B2(G472), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n359), .B1(new_n360), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n357), .A2(new_n629), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NOR2_X1   g487(.A1(new_n308), .A2(new_n312), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n668), .B(KEYINPUT39), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT96), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT38), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n600), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n642), .A2(new_n644), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n505), .B1(new_n491), .B2(new_n494), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n494), .A2(new_n505), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n294), .B1(new_n684), .B2(new_n517), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n515), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n357), .A2(new_n401), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n531), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n678), .A2(new_n679), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n215), .ZN(G45));
  NOR3_X1   g507(.A1(new_n666), .A2(new_n624), .A3(new_n668), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n665), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT97), .B(G146), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G48));
  NAND2_X1  g511(.A1(new_n303), .A2(new_n304), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n294), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(G469), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT98), .B1(new_n305), .B2(new_n187), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n300), .A2(new_n307), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n311), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n530), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n625), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n631), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  INV_X1    g525(.A(new_n531), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n598), .B2(new_n599), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n713), .A2(new_n311), .A3(new_n704), .A4(new_n703), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n666), .A2(new_n402), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n663), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT99), .B(G119), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G21));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n688), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n605), .A2(KEYINPUT100), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n604), .A2(new_n722), .A3(G472), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n500), .B(new_n508), .C1(new_n518), .C2(new_n498), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n510), .A3(new_n294), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n458), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n720), .A2(new_n705), .A3(new_n727), .A4(new_n363), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NOR2_X1   g543(.A1(new_n682), .A2(new_n726), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n624), .A2(new_n668), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n714), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  AOI21_X1  g547(.A(KEYINPUT101), .B1(new_n283), .B2(new_n287), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n293), .B2(KEYINPUT101), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n312), .B1(new_n736), .B2(new_n704), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n600), .A2(new_n712), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n530), .A4(new_n731), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT102), .B(G131), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G33));
  XNOR2_X1  g557(.A(new_n670), .B(KEYINPUT103), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n737), .A3(new_n530), .A4(new_n738), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  XNOR2_X1  g560(.A(new_n738), .B(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n620), .A2(new_n357), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT43), .Z(new_n749));
  INV_X1    g563(.A(new_n682), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n635), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n752), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n747), .B(KEYINPUT105), .C1(new_n751), .C2(new_n752), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n187), .B1(new_n293), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n704), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n311), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n675), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n755), .A2(new_n772), .A3(new_n756), .A4(new_n757), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n759), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n311), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n738), .A2(new_n731), .A3(new_n458), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n666), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  AND2_X1   g595(.A1(new_n703), .A2(new_n704), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n311), .A2(new_n531), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n687), .A2(new_n748), .A3(new_n458), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n783), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n681), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n397), .B2(new_n400), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n609), .A2(new_n365), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT107), .A3(new_n399), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n357), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n362), .B1(new_n624), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n607), .A2(new_n595), .A3(new_n601), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n635), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n642), .A2(new_n644), .A3(new_n636), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT94), .B1(new_n655), .B2(new_n656), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n402), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n674), .A2(new_n595), .A3(new_n601), .A4(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n602), .B(new_n797), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n659), .B(new_n403), .C1(new_n658), .C2(new_n530), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT108), .B1(new_n807), .B2(new_n797), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n530), .B(new_n705), .C1(new_n625), .C2(new_n631), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n716), .A2(new_n810), .A3(new_n728), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n730), .A2(new_n731), .A3(new_n738), .A4(new_n737), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n791), .A2(new_n669), .A3(new_n793), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n623), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n598), .A3(new_n531), .A4(new_n599), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n666), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n663), .A2(new_n674), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n818), .A3(new_n745), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n820), .A3(new_n741), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT109), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n739), .B(KEYINPUT42), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n811), .A3(new_n819), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n804), .A2(new_n805), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n807), .A2(KEYINPUT108), .A3(new_n797), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n663), .B(new_n664), .C1(new_n694), .C2(new_n671), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n736), .A2(new_n704), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n654), .A2(new_n312), .A3(new_n643), .A4(new_n668), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n720), .A2(new_n687), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n732), .A3(new_n833), .A4(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(new_n732), .A3(new_n833), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n822), .A2(new_n829), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT111), .B1(new_n838), .B2(KEYINPUT53), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n822), .A2(new_n829), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n839), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n838), .A2(KEYINPUT111), .A3(KEYINPUT53), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n789), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n749), .A2(new_n359), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n705), .A2(new_n738), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n530), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT48), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n714), .A3(new_n727), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(G952), .A3(new_n285), .ZN(new_n853));
  INV_X1    g667(.A(new_n359), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n687), .A2(new_n458), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n851), .B(new_n853), .C1(new_n624), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n727), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n681), .A2(new_n712), .A3(new_n705), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT50), .Z(new_n861));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n730), .A3(new_n849), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT112), .Z(new_n863));
  NOR3_X1   g677(.A1(new_n856), .A2(new_n623), .A3(new_n620), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n778), .B1(new_n312), .B2(new_n782), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n747), .A2(new_n848), .A3(new_n727), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n857), .B1(new_n869), .B2(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n868), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n871), .A2(KEYINPUT113), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT113), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n843), .A2(new_n842), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT53), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n838), .A2(KEYINPUT53), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n847), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n788), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n837), .A2(new_n834), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n828), .B1(new_n824), .B2(new_n827), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n887), .B2(new_n840), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n294), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n585), .A2(new_n588), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n587), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n892), .A2(new_n896), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n285), .A2(G952), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G51));
  XNOR2_X1  g714(.A(new_n888), .B(new_n789), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n764), .B(KEYINPUT57), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n698), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n763), .B(KEYINPUT115), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n889), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n899), .B1(new_n904), .B2(new_n906), .ZN(G54));
  AND2_X1   g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n878), .A2(G902), .A3(new_n347), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n899), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n841), .B2(new_n884), .ZN(new_n912));
  OAI211_X1 g726(.A(G902), .B(new_n908), .C1(new_n912), .C2(new_n883), .ZN(new_n913));
  INV_X1    g727(.A(new_n347), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(KEYINPUT116), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT116), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT117), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n911), .B(new_n919), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(G60));
  XOR2_X1   g735(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n922));
  NOR2_X1   g736(.A1(new_n364), .A2(new_n294), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n901), .A2(new_n617), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n910), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n847), .B2(new_n879), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n618), .ZN(G63));
  XNOR2_X1  g742(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT119), .Z(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n931), .B1(new_n888), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n455), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT120), .B(new_n934), .C1(new_n912), .C2(new_n883), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n910), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n639), .B1(new_n936), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n930), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n640), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n910), .A3(new_n939), .A4(new_n929), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(G66));
  INV_X1    g760(.A(G224), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n361), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n809), .A2(new_n811), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(G953), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n893), .B1(G898), .B2(new_n285), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT122), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n950), .B(new_n953), .ZN(G69));
  AOI21_X1  g768(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n480), .B1(new_n490), .B2(KEYINPUT30), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n327), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n774), .A2(new_n780), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n624), .A2(new_n795), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n738), .A2(new_n530), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n677), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n830), .A2(new_n732), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n692), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n692), .B2(new_n963), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n958), .B(new_n966), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n957), .B1(new_n970), .B2(new_n285), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n741), .A2(new_n745), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n719), .A2(new_n666), .A3(new_n458), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n962), .B(new_n976), .C1(new_n771), .C2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n958), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n774), .A2(new_n978), .A3(new_n780), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT126), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n285), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n957), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(G900), .B2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n971), .B2(new_n972), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n955), .B1(new_n974), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n971), .A2(new_n972), .ZN(new_n988));
  INV_X1    g802(.A(new_n955), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n973), .A3(new_n989), .A4(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  INV_X1    g807(.A(new_n949), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(new_n970), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n899), .B1(new_n995), .B2(new_n683), .ZN(new_n996));
  INV_X1    g810(.A(new_n993), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n979), .A2(new_n981), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(new_n949), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n491), .A2(new_n494), .A3(new_n505), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n499), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n993), .B1(new_n525), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT127), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n845), .B2(new_n846), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1001), .A2(new_n1005), .ZN(G57));
endmodule


