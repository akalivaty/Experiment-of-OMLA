//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929;
  NAND3_X1  g000(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT24), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n203), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT68), .B1(new_n212), .B2(new_n202), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT69), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT25), .B1(new_n215), .B2(KEYINPUT23), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n218), .A2(G169gat), .A3(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n220), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n216), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n212), .A2(new_n202), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n205), .A2(KEYINPUT24), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n204), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n203), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n204), .A2(new_n207), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(new_n202), .A3(new_n212), .ZN(new_n236));
  INV_X1    g035(.A(new_n215), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n221), .B1(new_n237), .B2(new_n218), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n215), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n236), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n210), .A2(KEYINPUT27), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(new_n211), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT27), .B(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n211), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n249), .A2(new_n252), .A3(new_n204), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n220), .B1(new_n215), .B2(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n255), .A2(KEYINPUT70), .B1(new_n254), .B2(new_n215), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(KEYINPUT70), .B2(new_n255), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n244), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G113gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n263), .A3(G120gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n260), .A2(G120gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G134gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  INV_X1    g073(.A(G120gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G113gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n267), .A2(new_n273), .B1(new_n277), .B2(new_n272), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n234), .A2(new_n243), .B1(new_n257), .B2(new_n253), .ZN(new_n281));
  INV_X1    g080(.A(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT32), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G15gat), .B(G43gat), .Z(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(KEYINPUT32), .C1(new_n286), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n280), .B1(new_n279), .B2(new_n283), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n295), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(new_n291), .A3(new_n293), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT36), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n298), .A3(new_n301), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n294), .A2(KEYINPUT73), .A3(new_n297), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(KEYINPUT36), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT0), .ZN(new_n309));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G141gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT81), .B1(new_n312), .B2(G148gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(new_n316), .A3(KEYINPUT82), .A4(new_n317), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(KEYINPUT79), .B2(KEYINPUT2), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n315), .A2(G141gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n312), .A2(G148gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n329), .A2(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(KEYINPUT78), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(G155gat), .A3(G162gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n336), .A2(new_n338), .B1(new_n323), .B2(new_n324), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n334), .B2(new_n339), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n328), .B(new_n278), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n346), .A2(new_n322), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n315), .A2(G141gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n330), .B1(new_n317), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n336), .A2(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n323), .A2(new_n324), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT80), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n328), .A4(new_n278), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n344), .A2(new_n345), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n328), .B1(new_n340), .B2(new_n341), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(KEYINPUT83), .A3(new_n328), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT3), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n318), .A2(new_n319), .B1(new_n326), .B2(new_n325), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n353), .A2(new_n354), .B1(new_n321), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n278), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n357), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(new_n361), .A3(new_n282), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n345), .B1(new_n369), .B2(new_n342), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n357), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n368), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(KEYINPUT6), .B(new_n311), .C1(new_n371), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377));
  INV_X1    g176(.A(new_n311), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n371), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n373), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n369), .A2(new_n342), .ZN(new_n382));
  INV_X1    g181(.A(new_n345), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n368), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n378), .B1(new_n386), .B2(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n376), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G197gat), .B(G204gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT22), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n391), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G226gat), .ZN(new_n399));
  INV_X1    g198(.A(G233gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n259), .A2(KEYINPUT75), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT75), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n281), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n281), .B2(KEYINPUT29), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n398), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n259), .A2(new_n401), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n413), .A3(new_n398), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n408), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n388), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT76), .B1(new_n408), .B2(new_n415), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n259), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n402), .A2(new_n405), .B1(new_n424), .B2(new_n404), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n422), .B(new_n414), .C1(new_n425), .C2(new_n398), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n412), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(KEYINPUT30), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT77), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT77), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n364), .A2(new_n365), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n398), .B1(new_n432), .B2(new_n423), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n360), .A2(new_n361), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n365), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G228gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n396), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(new_n389), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT29), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n392), .A2(KEYINPUT86), .A3(new_n395), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n389), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT3), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n437), .B1(new_n444), .B2(new_n364), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n436), .A2(new_n437), .B1(new_n433), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(G22gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(G22gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449));
  INV_X1    g248(.A(G50gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT87), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n448), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n446), .A2(G22gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n307), .B1(new_n431), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n380), .B2(new_n387), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n311), .B1(new_n371), .B2(new_n375), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n311), .B1(new_n367), .B2(new_n368), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT6), .B1(new_n467), .B2(new_n386), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT88), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n416), .B1(new_n387), .B2(KEYINPUT6), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(new_n414), .C1(new_n425), .C2(new_n398), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n407), .A2(new_n413), .A3(new_n397), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT37), .B(new_n473), .C1(new_n425), .C2(new_n397), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n412), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n465), .A2(new_n469), .A3(new_n470), .A4(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n476), .A2(new_n376), .A3(new_n417), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(KEYINPUT89), .A3(new_n465), .A4(new_n469), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n421), .A2(KEYINPUT37), .A3(new_n426), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n472), .A2(new_n412), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT38), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT90), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT38), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n479), .A2(new_n481), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n461), .A2(new_n456), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n344), .A2(new_n356), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n345), .B1(new_n373), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT39), .B1(new_n382), .B2(new_n383), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n494), .B(new_n378), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n498), .A2(new_n499), .A3(new_n387), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n419), .A2(new_n427), .A3(new_n428), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n463), .B1(new_n489), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n490), .A2(new_n306), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n431), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n298), .A2(new_n301), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n462), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(new_n501), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n465), .A2(new_n469), .A3(new_n376), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n505), .A2(KEYINPUT35), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G43gat), .B(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT92), .ZN(new_n516));
  OR3_X1    g315(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n519), .B(new_n520), .C1(KEYINPUT15), .C2(new_n514), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n523), .A2(new_n524), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n516), .A2(new_n521), .B1(new_n525), .B2(new_n515), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n527), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT93), .Z(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n532), .B2(new_n526), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT13), .Z(new_n537));
  AND2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n526), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n532), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n536), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT12), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n553), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  AOI21_X1  g366(.A(new_n532), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT97), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n576), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n582), .A2(new_n591), .A3(new_n583), .A4(new_n587), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n541), .A2(new_n543), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n595), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT101), .B1(new_n598), .B2(new_n600), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT98), .ZN(new_n606));
  XOR2_X1   g405(.A(G134gat), .B(G162gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n598), .A2(new_n600), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n603), .A2(new_n604), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n601), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n579), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G230gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n400), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n593), .B(new_n564), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n564), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n618), .A2(new_n616), .A3(new_n400), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n557), .A2(new_n615), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n513), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n388), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n501), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G8gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(G8gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n634), .A2(new_n646), .A3(new_n506), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n513), .A2(new_n307), .A3(new_n633), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n490), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT103), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT43), .B(G22gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n614), .B1(new_n503), .B2(new_n512), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n489), .A2(new_n502), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n431), .B2(new_n462), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(KEYINPUT105), .A3(new_n490), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n656), .A2(new_n307), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n508), .A2(new_n511), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n614), .B(KEYINPUT106), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT44), .ZN(new_n668));
  AOI22_X1  g467(.A1(KEYINPUT44), .A2(new_n655), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n557), .ZN(new_n670));
  INV_X1    g469(.A(new_n579), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n670), .A2(new_n671), .A3(new_n631), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n654), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n614), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n490), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n656), .A2(new_n676), .A3(new_n307), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(new_n664), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n668), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n661), .B2(new_n664), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT107), .B(new_n672), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n388), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n678), .A2(new_n672), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n388), .A2(G29gat), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT104), .B1(new_n686), .B2(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(KEYINPUT45), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n685), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n685), .A2(KEYINPUT108), .A3(new_n690), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1328gat));
  INV_X1    g497(.A(new_n501), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n684), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n686), .A2(G36gat), .A3(new_n699), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n669), .A2(new_n673), .ZN(new_n705));
  INV_X1    g504(.A(new_n307), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  AOI211_X1 g507(.A(G43gat), .B(new_n686), .C1(new_n301), .C2(new_n298), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n674), .A2(new_n706), .A3(new_n683), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n711), .A2(KEYINPUT109), .A3(G43gat), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n711), .B2(G43gat), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n709), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g514(.A1(new_n686), .A2(G50gat), .A3(new_n462), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n674), .A2(new_n490), .A3(new_n683), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(G50gat), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n450), .B1(new_n705), .B2(new_n490), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n718), .A2(KEYINPUT48), .B1(new_n719), .B2(new_n721), .ZN(G1331gat));
  NAND3_X1  g521(.A1(new_n670), .A2(new_n615), .A3(new_n631), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT110), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n665), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n727), .A3(new_n665), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n635), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g530(.A(new_n699), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n726), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT112), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT112), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n729), .A2(new_n741), .A3(new_n506), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n728), .ZN(new_n743));
  OAI21_X1  g542(.A(G71gat), .B1(new_n743), .B2(new_n307), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n490), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n670), .A2(new_n579), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT113), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n614), .A3(new_n665), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n631), .A2(new_n635), .A3(new_n585), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n751), .A2(new_n631), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n669), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n585), .B1(new_n760), .B2(new_n635), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n757), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n757), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1336gat));
  NOR3_X1   g563(.A1(new_n632), .A2(new_n699), .A3(G92gat), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n759), .A2(new_n669), .A3(new_n699), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n586), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT52), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n586), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(G1337gat));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n631), .A2(new_n775), .A3(new_n506), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT116), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n754), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n759), .A2(new_n669), .A3(new_n307), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n775), .B2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n632), .A2(G106gat), .A3(new_n462), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n754), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n760), .B2(new_n490), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT53), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1339gat));
  NAND4_X1  g586(.A1(new_n615), .A2(new_n554), .A3(new_n556), .A4(new_n632), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n545), .A2(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n552), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n556), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n627), .B1(new_n622), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n622), .A2(new_n796), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n620), .A2(new_n621), .A3(new_n617), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n629), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(new_n666), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n557), .A2(new_n803), .B1(new_n795), .B2(new_n631), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n666), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n790), .B1(new_n806), .B2(new_n579), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n388), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n504), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n699), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n261), .A3(new_n263), .A4(new_n557), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n508), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n670), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1340gat));
  NAND2_X1  g613(.A1(new_n631), .A2(new_n275), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT119), .Z(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G120gat), .B1(new_n812), .B2(new_n632), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  NAND3_X1  g618(.A1(new_n810), .A2(new_n270), .A3(new_n671), .ZN(new_n820));
  OAI21_X1  g619(.A(G127gat), .B1(new_n812), .B2(new_n579), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1342gat));
  NAND2_X1  g621(.A1(new_n699), .A2(new_n614), .ZN(new_n823));
  AOI211_X1 g622(.A(G134gat), .B(new_n823), .C1(KEYINPUT120), .C2(KEYINPUT56), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n812), .B2(new_n675), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(KEYINPUT121), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(KEYINPUT121), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n827), .B(new_n828), .C1(new_n830), .C2(new_n831), .ZN(G1343gat));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n806), .A2(new_n579), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n833), .B(new_n490), .C1(new_n834), .C2(new_n790), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n804), .B1(new_n805), .B2(new_n614), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n790), .B1(new_n836), .B2(new_n579), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n462), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n706), .A2(new_n388), .A3(new_n501), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G141gat), .B1(new_n840), .B2(new_n670), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n706), .A2(new_n462), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n808), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n501), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n670), .A2(G141gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(KEYINPUT122), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(KEYINPUT58), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n841), .B(new_n846), .C1(KEYINPUT122), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n315), .A2(KEYINPUT59), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n844), .B2(new_n631), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n840), .A2(new_n632), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n805), .A2(new_n614), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n795), .A2(new_n614), .A3(new_n803), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n671), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n788), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n833), .B(new_n490), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n807), .B2(new_n462), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n631), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n839), .A2(KEYINPUT59), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n855), .A2(KEYINPUT59), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n854), .B1(new_n864), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g664(.A(G155gat), .B1(new_n840), .B2(new_n579), .ZN(new_n866));
  INV_X1    g665(.A(new_n844), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n671), .A2(new_n323), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n866), .B(KEYINPUT123), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1346gat));
  NOR3_X1   g672(.A1(new_n843), .A2(G162gat), .A3(new_n823), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT124), .ZN(new_n875));
  OAI21_X1  g674(.A(G162gat), .B1(new_n840), .B2(new_n667), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n699), .A2(new_n635), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n807), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n504), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n557), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n807), .A2(new_n507), .A3(new_n879), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n557), .A2(G169gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1348gat));
  NOR3_X1   g685(.A1(new_n881), .A2(G176gat), .A3(new_n632), .ZN(new_n887));
  INV_X1    g686(.A(G176gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n884), .B2(new_n631), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n887), .A2(new_n889), .ZN(G1349gat));
  AND4_X1   g689(.A1(new_n250), .A2(new_n880), .A3(new_n504), .A4(new_n671), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n210), .B1(new_n884), .B2(new_n671), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n211), .A3(new_n666), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n211), .B1(new_n884), .B2(new_n614), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1351gat));
  NOR2_X1   g699(.A1(new_n706), .A2(new_n879), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n860), .A2(new_n861), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G197gat), .B1(new_n902), .B2(new_n670), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n807), .A2(new_n462), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n670), .A2(G197gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n904), .A2(KEYINPUT126), .A3(new_n901), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n904), .A2(new_n901), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(G204gat), .A3(new_n632), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  INV_X1    g717(.A(new_n901), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n862), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1353gat));
  OR3_X1    g720(.A1(new_n916), .A2(G211gat), .A3(new_n579), .ZN(new_n922));
  OAI21_X1  g721(.A(G211gat), .B1(new_n902), .B2(new_n579), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1354gat));
  OAI21_X1  g726(.A(G218gat), .B1(new_n902), .B2(new_n675), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n667), .A2(G218gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n916), .B2(new_n929), .ZN(G1355gat));
endmodule


