//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  OR2_X1    g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(new_n203), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n205), .C1(new_n208), .C2(KEYINPUT2), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n215));
  XNOR2_X1  g014(.A(G197gat), .B(G204gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G197gat), .B(G204gat), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT73), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n218), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n222), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT75), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n225), .B1(new_n230), .B2(new_n215), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n229), .A2(new_n218), .B1(new_n231), .B2(new_n224), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n214), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT85), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n227), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n243), .B2(new_n213), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n244), .B2(new_n210), .ZN(new_n245));
  NAND2_X1  g044(.A1(G228gat), .A2(G233gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n215), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n229), .B2(new_n218), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n233), .B1(new_n225), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n250), .B2(new_n213), .ZN(new_n251));
  OAI211_X1 g050(.A(G228gat), .B(G233gat), .C1(new_n251), .C2(new_n210), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n237), .B1(new_n221), .B2(new_n226), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT75), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n236), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(new_n255), .B1(new_n213), .B2(new_n212), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n252), .A2(new_n256), .A3(KEYINPUT86), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n211), .B1(new_n253), .B2(KEYINPUT29), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n207), .A2(new_n209), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n246), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n239), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n247), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G22gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT31), .B(G50gat), .Z(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G22gat), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n247), .B(new_n269), .C1(new_n257), .C2(new_n262), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n270), .B2(KEYINPUT88), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT87), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT86), .B1(new_n252), .B2(new_n256), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n261), .A2(new_n258), .A3(new_n239), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n274), .A2(new_n275), .B1(new_n246), .B2(new_n245), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n273), .B1(new_n276), .B2(new_n269), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n265), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n272), .A3(new_n268), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n276), .B2(new_n269), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n264), .C1(new_n281), .C2(new_n268), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT32), .ZN(new_n284));
  OR3_X1    g083(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(G169gat), .ZN(new_n287));
  INV_X1    g086(.A(G176gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT65), .B(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT27), .B1(new_n295), .B2(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n291), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n302), .B(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n311), .C1(new_n287), .C2(new_n288), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n304), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n290), .A2(new_n295), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n314), .B(KEYINPUT25), .C1(new_n315), .C2(new_n306), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(G113gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n327), .A2(new_n328), .B1(KEYINPUT67), .B2(new_n319), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(G113gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n320), .A2(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n319), .A2(KEYINPUT67), .ZN(new_n334));
  INV_X1    g133(.A(new_n328), .ZN(new_n335));
  NOR2_X1   g134(.A1(G127gat), .A2(G134gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n338), .A3(KEYINPUT68), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n318), .A2(KEYINPUT69), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n302), .A2(new_n301), .B1(new_n313), .B2(new_n316), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n339), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n284), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n350), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT70), .ZN(new_n357));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G43gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT72), .B(G15gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n354), .A2(new_n363), .A3(new_n355), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n353), .A2(new_n357), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n351), .B1(new_n355), .B2(new_n361), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n349), .A2(new_n350), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(KEYINPUT34), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n365), .A3(new_n366), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n283), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374));
  AND2_X1   g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n318), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n345), .A2(KEYINPUT29), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n375), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n234), .A2(new_n238), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n376), .C1(new_n377), .C2(new_n375), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n381), .B2(new_n382), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n382), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n391), .A2(KEYINPUT30), .A3(new_n385), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n374), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n388), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT89), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT76), .B1(new_n210), .B2(new_n211), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n330), .A2(new_n338), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n260), .A2(new_n404), .A3(KEYINPUT3), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n212), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n403), .A2(new_n410), .A3(new_n260), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT77), .B1(new_n210), .B2(new_n340), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT4), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n346), .A2(new_n414), .A3(new_n210), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  AOI211_X1 g216(.A(KEYINPUT4), .B(new_n260), .C1(new_n342), .C2(new_n339), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(KEYINPUT81), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n410), .B1(new_n403), .B2(new_n260), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n210), .A2(KEYINPUT77), .A3(new_n340), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT81), .B1(new_n423), .B2(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n415), .A2(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT82), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n401), .B(new_n408), .C1(new_n420), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n411), .A2(new_n412), .B1(new_n340), .B2(new_n210), .ZN(new_n434));
  INV_X1    g233(.A(new_n407), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT79), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT5), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT78), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n414), .B1(new_n411), .B2(new_n412), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n408), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n442), .A2(new_n407), .A3(new_n406), .A4(new_n443), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT78), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n438), .A2(new_n440), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n427), .A2(new_n433), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n433), .B1(new_n427), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n400), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n427), .A2(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n432), .ZN(new_n453));
  INV_X1    g252(.A(new_n400), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n373), .A2(new_n399), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n283), .A2(new_n371), .A3(new_n372), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n396), .A2(new_n397), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n455), .A4(new_n459), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n457), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n278), .A2(new_n282), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n381), .A2(new_n469), .A3(new_n382), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n470), .A2(new_n385), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n391), .A2(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n450), .B2(new_n455), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n381), .A2(KEYINPUT90), .A3(new_n382), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(KEYINPUT37), .C1(KEYINPUT90), .C2(new_n381), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n471), .A3(new_n468), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n477), .A2(new_n395), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n467), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n434), .A2(new_n435), .ZN(new_n480));
  INV_X1    g279(.A(new_n406), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n417), .B1(new_n416), .B2(new_n419), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n424), .A2(KEYINPUT82), .A3(new_n425), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT39), .B(new_n480), .C1(new_n484), .C2(new_n407), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n406), .B1(new_n420), .B2(new_n426), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n435), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n433), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n449), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n485), .A2(KEYINPUT40), .A3(new_n488), .A4(new_n433), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n399), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n466), .B1(new_n479), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n473), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n427), .A2(new_n433), .A3(new_n447), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n454), .B1(new_n453), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n449), .A2(new_n400), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n478), .B(new_n495), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n466), .A2(new_n493), .A3(new_n499), .A4(new_n283), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n462), .A2(new_n463), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(new_n371), .ZN(new_n504));
  INV_X1    g303(.A(new_n372), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n371), .A2(KEYINPUT36), .A3(new_n372), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n502), .A2(new_n467), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n465), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT16), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n510), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT100), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(G64gat), .ZN(new_n520));
  INV_X1    g319(.A(G64gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(G57gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(G57gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(G64gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT100), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT101), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n520), .B2(new_n522), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n529), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT101), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n516), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n295), .ZN(new_n541));
  INV_X1    g340(.A(G231gat), .ZN(new_n542));
  INV_X1    g341(.A(G233gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n540), .B(G183gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G127gat), .B(G155gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT20), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n549), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n539), .A2(new_n517), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G211gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n554), .B(new_n556), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n553), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  INV_X1    g358(.A(G36gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT14), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT14), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G50gat), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT15), .B1(new_n566), .B2(G43gat), .ZN(new_n567));
  INV_X1    g366(.A(G43gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G50gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(KEYINPUT94), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G43gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n574), .A3(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(G50gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n577), .A2(new_n578), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n562), .A2(G29gat), .A3(G36gat), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT14), .B1(new_n559), .B2(new_n560), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT95), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n570), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n571), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(G99gat), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT8), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n589), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n593), .B(KEYINPUT7), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(new_n597), .A3(new_n589), .A4(new_n592), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n588), .A2(new_n603), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n579), .A2(new_n585), .ZN(new_n607));
  INV_X1    g406(.A(new_n571), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n587), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI211_X1 g408(.A(KEYINPUT96), .B(new_n571), .C1(new_n579), .C2(new_n585), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n586), .A2(KEYINPUT17), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n602), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(KEYINPUT103), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n605), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(KEYINPUT103), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n623), .A3(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n509), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n630));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n516), .A3(new_n612), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n516), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n588), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n635), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n637), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n588), .A2(new_n638), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n588), .A2(new_n638), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n636), .A2(KEYINPUT18), .A3(new_n639), .A4(new_n637), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n644), .A2(new_n651), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT100), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT100), .B1(new_n524), .B2(new_n525), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n530), .B1(new_n657), .B2(KEYINPUT9), .ZN(new_n658));
  INV_X1    g457(.A(new_n538), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n602), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n532), .A2(new_n601), .A3(new_n599), .A4(new_n538), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n527), .B2(new_n531), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n603), .A3(new_n665), .A4(KEYINPUT10), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n662), .B2(new_n661), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n660), .A2(new_n662), .ZN(new_n671));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n654), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n629), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n450), .A2(new_n455), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n511), .ZN(G1324gat));
  INV_X1    g489(.A(new_n399), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n693));
  OR2_X1    g492(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n697), .B(new_n698), .C1(new_n515), .C2(new_n692), .ZN(G1325gat));
  INV_X1    g498(.A(new_n683), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n504), .A2(new_n505), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n506), .A2(new_n507), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT106), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT107), .Z(new_n706));
  AOI21_X1  g505(.A(new_n702), .B1(new_n700), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n683), .A2(new_n283), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NAND3_X1  g509(.A1(new_n493), .A2(new_n499), .A3(new_n283), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT91), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n502), .A2(new_n467), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n493), .A2(new_n499), .A3(new_n466), .A4(new_n283), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n703), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n716));
  INV_X1    g515(.A(new_n457), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n627), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n558), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n682), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n559), .A3(new_n687), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n509), .B2(new_n627), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n719), .A2(KEYINPUT44), .A3(new_n720), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n723), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n732), .B2(new_n688), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n726), .A2(new_n733), .ZN(G1328gat));
  NAND3_X1  g533(.A1(new_n724), .A2(new_n560), .A3(new_n399), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n732), .B2(new_n691), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1329gat));
  AND2_X1   g538(.A1(new_n572), .A2(new_n574), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n732), .B2(new_n703), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n742), .A3(new_n701), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n743), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n704), .A3(new_n731), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n740), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(KEYINPUT47), .B2(new_n747), .ZN(G1330gat));
  NAND2_X1  g547(.A1(new_n467), .A2(G50gat), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n721), .A2(new_n283), .A3(new_n723), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n732), .A2(new_n749), .B1(G50gat), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g551(.A(new_n654), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n628), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n719), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n681), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n687), .B(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n691), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  INV_X1    g564(.A(G71gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n704), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n756), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n757), .A2(new_n701), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1334gat));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n283), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT111), .B(G78gat), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n558), .A2(new_n753), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n728), .A2(new_n681), .A3(new_n729), .A4(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(G85gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n688), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n719), .A2(new_n720), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n719), .A2(new_n782), .A3(new_n720), .A4(new_n776), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n681), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n687), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n779), .B1(new_n785), .B2(new_n778), .ZN(G1336gat));
  OAI21_X1  g585(.A(G92gat), .B1(new_n777), .B2(new_n691), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n691), .A2(G92gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n781), .A2(new_n681), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n787), .B(new_n791), .C1(new_n788), .C2(KEYINPUT52), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n784), .A2(new_n590), .A3(new_n701), .ZN(new_n796));
  OAI21_X1  g595(.A(G99gat), .B1(new_n777), .B2(new_n767), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n784), .A2(new_n591), .A3(new_n467), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G106gat), .B1(new_n777), .B2(new_n283), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT53), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n799), .B(new_n802), .C1(new_n800), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1339gat));
  NAND4_X1  g606(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n672), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n668), .A2(new_n810), .A3(new_n669), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n677), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n680), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n668), .A2(new_n669), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(KEYINPUT54), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n677), .B(new_n811), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n816), .A2(KEYINPUT114), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT114), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n653), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n644), .A2(new_n651), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n642), .A2(new_n635), .A3(new_n649), .A4(new_n650), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n647), .A2(new_n648), .A3(new_n646), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n637), .B1(new_n636), .B2(new_n639), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n634), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n681), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n824), .A2(new_n830), .A3(new_n827), .A4(new_n681), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n627), .B1(new_n823), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n824), .A2(new_n827), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n625), .A3(new_n626), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n820), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n558), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n628), .A2(new_n753), .A3(new_n681), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n373), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n691), .A3(new_n758), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n320), .A3(new_n753), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n688), .A2(new_n399), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n320), .B1(new_n847), .B2(new_n753), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  INV_X1    g650(.A(new_n681), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n681), .A2(new_n322), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n842), .B2(new_n854), .ZN(G1341gat));
  NOR3_X1   g654(.A1(new_n846), .A2(new_n325), .A3(new_n722), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n843), .A2(new_n558), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n325), .ZN(G1342gat));
  NOR3_X1   g657(.A1(new_n842), .A2(G134gat), .A3(new_n627), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n846), .B2(new_n627), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n816), .A2(new_n817), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n813), .B(new_n864), .C1(new_n652), .C2(new_n653), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n828), .A2(KEYINPUT117), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n834), .A2(new_n867), .A3(new_n681), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n836), .B1(new_n869), .B2(new_n627), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n863), .B1(new_n870), .B2(new_n558), .ZN(new_n871));
  INV_X1    g670(.A(new_n839), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n828), .B(new_n867), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n720), .B1(new_n873), .B2(new_n865), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT118), .B(new_n722), .C1(new_n874), .C2(new_n836), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n283), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n467), .B1(new_n838), .B2(new_n839), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n845), .A2(new_n703), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT119), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n876), .A2(new_n878), .B1(new_n880), .B2(new_n877), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n753), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(G141gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n882), .A2(KEYINPUT119), .A3(new_n884), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n886), .B2(new_n883), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n654), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(G141gat), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT120), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n840), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n758), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n399), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n283), .B(new_n704), .C1(new_n898), .C2(KEYINPUT121), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n895), .A4(new_n753), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n891), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n886), .A2(new_n654), .A3(new_n883), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n902), .B(new_n905), .C1(new_n895), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(G1344gat));
  AND2_X1   g707(.A1(new_n900), .A2(new_n901), .ZN(new_n909));
  INV_X1    g708(.A(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n681), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n839), .B(KEYINPUT122), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n870), .A2(new_n558), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n877), .B(new_n467), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n681), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(new_n883), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n852), .B1(new_n892), .B2(new_n893), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(KEYINPUT59), .A3(new_n910), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n911), .B1(new_n919), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(G155gat), .B1(new_n909), .B2(new_n558), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n722), .B1(new_n892), .B2(new_n893), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(G155gat), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(new_n720), .B1(new_n885), .B2(new_n888), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(G162gat), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G162gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n931), .A3(new_n720), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n758), .A2(new_n691), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n841), .ZN(new_n935));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n654), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n840), .A2(new_n687), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n458), .A2(new_n399), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT124), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n938), .A2(KEYINPUT124), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n287), .A3(new_n753), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n936), .A2(new_n943), .ZN(G1348gat));
  NOR3_X1   g743(.A1(new_n935), .A2(new_n288), .A3(new_n852), .ZN(new_n945));
  AOI21_X1  g744(.A(G176gat), .B1(new_n942), .B2(new_n681), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n935), .B2(new_n722), .ZN(new_n948));
  INV_X1    g747(.A(new_n299), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n941), .A2(new_n722), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n720), .A3(new_n290), .ZN(new_n956));
  OAI21_X1  g755(.A(G190gat), .B1(new_n935), .B2(new_n627), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  AND4_X1   g759(.A1(new_n467), .A2(new_n937), .A3(new_n399), .A4(new_n767), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  INV_X1    g761(.A(G197gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n963), .A3(new_n753), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n704), .A2(new_n691), .A3(new_n758), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n915), .A3(new_n916), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n966), .A2(KEYINPUT127), .A3(new_n654), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(new_n966), .B2(new_n654), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(G197gat), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n964), .A2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n961), .A2(new_n971), .A3(new_n681), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  INV_X1    g772(.A(new_n965), .ZN(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n917), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1353gat));
  INV_X1    g775(.A(G211gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n977), .A3(new_n558), .ZN(new_n978));
  OAI21_X1  g777(.A(G211gat), .B1(new_n966), .B2(new_n722), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT63), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n962), .A2(new_n984), .A3(new_n720), .ZN(new_n985));
  OAI21_X1  g784(.A(G218gat), .B1(new_n966), .B2(new_n627), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


