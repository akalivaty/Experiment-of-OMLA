//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n190), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G134), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT11), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n201), .A3(G134), .ZN(new_n206));
  AOI211_X1 g020(.A(G131), .B(new_n202), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n206), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(G137), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT0), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(KEYINPUT0), .B2(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT65), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n221), .B2(G146), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(G143), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n228), .A2(new_n226), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n220), .A2(new_n227), .B1(new_n229), .B2(new_n216), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n200), .B1(new_n213), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n201), .B2(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n201), .A2(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n210), .A2(new_n240), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n209), .A2(new_n208), .A3(new_n210), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT70), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT28), .B1(new_n231), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n220), .A2(new_n227), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n229), .A2(new_n216), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n212), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n200), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n230), .B(new_n256), .C1(new_n207), .C2(new_n211), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n249), .A2(new_n254), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n245), .A2(new_n246), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n235), .A2(new_n228), .A3(new_n226), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n233), .B2(new_n227), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n212), .A2(new_n253), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n200), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n250), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT71), .B(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(G210), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT30), .A4(new_n257), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n200), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n272), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n250), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n249), .A2(new_n254), .A3(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n200), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n258), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT75), .B1(new_n285), .B2(KEYINPUT28), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n287), .B(new_n288), .C1(new_n284), .C2(new_n258), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n282), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G472), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n294), .B(KEYINPUT74), .Z(new_n295));
  NAND3_X1  g109(.A1(new_n278), .A2(new_n258), .A3(new_n273), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n278), .A2(new_n273), .A3(new_n298), .A4(new_n258), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(KEYINPUT31), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n288), .B1(new_n258), .B2(new_n263), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n272), .B1(new_n301), .B2(new_n250), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n278), .A2(new_n273), .A3(new_n303), .A4(new_n258), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI211_X1 g119(.A(KEYINPUT32), .B(new_n295), .C1(new_n300), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n305), .ZN(new_n308));
  INV_X1    g122(.A(new_n295), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n293), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(G234), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n319), .B1(new_n323), .B2(new_n317), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n224), .ZN(new_n325));
  OAI211_X1 g139(.A(G146), .B(new_n319), .C1(new_n323), .C2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n331), .A3(new_n335), .A4(new_n332), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G110), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT24), .B(G110), .Z(new_n338));
  XNOR2_X1  g152(.A(G119), .B(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n333), .A2(G110), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n326), .C1(G146), .C2(new_n323), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT77), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n347), .B1(new_n341), .B2(new_n343), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n314), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n343), .ZN(new_n354));
  INV_X1    g168(.A(new_n347), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n348), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n314), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n316), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n315), .A2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n312), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT25), .B1(new_n357), .B2(new_n314), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n352), .B(G902), .C1(new_n356), .C2(new_n348), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n315), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT78), .A3(new_n361), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n311), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n221), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n215), .A2(G143), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n203), .ZN(new_n375));
  INV_X1    g189(.A(G116), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT14), .A3(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(G116), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(G107), .B(new_n377), .C1(new_n379), .C2(KEYINPUT14), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n375), .B(new_n380), .C1(G107), .C2(new_n379), .ZN(new_n381));
  INV_X1    g195(.A(new_n372), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n382), .A2(KEYINPUT13), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n373), .B1(new_n382), .B2(KEYINPUT13), .ZN(new_n384));
  OAI21_X1  g198(.A(G134), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n374), .A2(new_n203), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n378), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n391), .A2(new_n313), .A3(G953), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(new_n314), .ZN(new_n394));
  INV_X1    g208(.A(G478), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(KEYINPUT15), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n314), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT15), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G478), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n267), .A2(G952), .ZN(new_n401));
  INV_X1    g215(.A(G234), .ZN(new_n402));
  INV_X1    g216(.A(G237), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n314), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT93), .B(G475), .Z(new_n411));
  XNOR2_X1  g225(.A(G113), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(G104), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(KEYINPUT71), .A2(G237), .ZN(new_n415));
  NOR2_X1   g229(.A1(KEYINPUT71), .A2(G237), .ZN(new_n416));
  OAI211_X1 g230(.A(G214), .B(new_n267), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT88), .B(G143), .Z(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n266), .A2(G214), .A3(new_n267), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT18), .A2(G131), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT89), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT90), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n419), .A2(new_n421), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n323), .B(new_n224), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n208), .B1(new_n419), .B2(new_n421), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(KEYINPUT91), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n327), .B1(KEYINPUT17), .B2(new_n430), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n419), .A2(new_n421), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(G131), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n439), .B2(KEYINPUT17), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n414), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n428), .A2(KEYINPUT91), .A3(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT91), .B1(new_n428), .B2(new_n431), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n414), .B(new_n440), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n436), .A2(KEYINPUT92), .A3(new_n414), .A4(new_n440), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n411), .B1(new_n448), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n323), .B(KEYINPUT19), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n439), .B(new_n326), .C1(G146), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n414), .B1(new_n436), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(G475), .A2(G902), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n446), .B2(new_n447), .ZN(new_n459));
  INV_X1    g273(.A(new_n457), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n449), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT94), .B(new_n449), .C1(new_n458), .C2(new_n461), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n410), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT3), .B1(new_n413), .B2(G107), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n387), .A3(G104), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n413), .A2(G107), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G101), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT80), .B(G101), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT4), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n476), .A3(G101), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n200), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n413), .A2(G107), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n387), .A2(G104), .ZN(new_n480));
  OAI21_X1  g294(.A(G101), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n376), .A2(G119), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT5), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n189), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(KEYINPUT82), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT82), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n329), .A2(G116), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n376), .A2(G119), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT5), .ZN(new_n491));
  OAI21_X1  g305(.A(G113), .B1(new_n489), .B2(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n482), .A2(new_n199), .A3(new_n487), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(G110), .B(G122), .Z(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT83), .ZN(new_n498));
  INV_X1    g312(.A(new_n496), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n478), .B2(new_n494), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n478), .A2(new_n494), .A3(new_n499), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT6), .ZN(new_n505));
  AND4_X1   g319(.A1(KEYINPUT84), .A2(new_n495), .A3(new_n505), .A4(new_n496), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT84), .B1(new_n500), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT86), .B1(new_n237), .B2(G125), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n261), .A2(new_n510), .A3(new_n321), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n253), .A2(G125), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  OR3_X1    g328(.A1(new_n230), .A2(KEYINPUT85), .A3(new_n321), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(G224), .A3(new_n267), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n267), .A2(G224), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n512), .A2(new_n514), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n508), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n496), .B(KEYINPUT8), .Z(new_n523));
  AOI22_X1  g337(.A1(new_n198), .A2(new_n195), .B1(new_n483), .B2(new_n486), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n474), .A2(new_n481), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND4_X1   g340(.A1(new_n199), .A2(new_n525), .A3(new_n493), .A4(new_n487), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n503), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n526), .A2(new_n527), .A3(new_n522), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n512), .B2(new_n513), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n533), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G210), .B1(G237), .B2(G902), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n521), .A2(new_n537), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  OAI21_X1  g358(.A(G221), .B1(new_n391), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(G469), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n525), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n239), .A2(new_n548), .A3(new_n248), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n232), .A2(G128), .B1(new_n228), .B2(new_n226), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n474), .B(new_n481), .C1(new_n550), .C2(new_n260), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n547), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n475), .A2(new_n230), .A3(new_n477), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n212), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G140), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n267), .A2(G227), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT81), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n261), .A2(new_n525), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n261), .B2(new_n525), .ZN(new_n563));
  INV_X1    g377(.A(new_n551), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n560), .B1(new_n565), .B2(new_n212), .ZN(new_n566));
  INV_X1    g380(.A(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n261), .A2(new_n525), .A3(new_n561), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n551), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n559), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n239), .A2(new_n548), .A3(new_n248), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n553), .A2(new_n552), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n213), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n558), .B1(new_n574), .B2(new_n554), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n546), .B(new_n314), .C1(new_n571), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n559), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(new_n554), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n566), .B2(new_n570), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n557), .B(KEYINPUT79), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n578), .B(G469), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n546), .A2(new_n314), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n576), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n371), .A2(new_n466), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(new_n473), .Z(G3));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n545), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n368), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n308), .A2(new_n309), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n308), .A2(new_n594), .A3(new_n314), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n300), .B2(new_n305), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n594), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n592), .B(new_n593), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n390), .A2(new_n392), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n601), .B2(KEYINPUT96), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(new_n393), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n603), .A2(KEYINPUT97), .A3(new_n395), .A4(G902), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT97), .B1(new_n394), .B2(G478), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n602), .B(new_n393), .Z(new_n606));
  NOR2_X1   g420(.A1(new_n395), .A2(G902), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n408), .ZN(new_n610));
  INV_X1    g424(.A(new_n542), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n539), .B1(new_n521), .B2(new_n537), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n610), .B(new_n544), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n464), .A2(new_n465), .A3(new_n609), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n600), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND3_X1  g435(.A1(new_n456), .A2(new_n450), .A3(new_n457), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT20), .B1(new_n459), .B2(new_n460), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n449), .A3(new_n400), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n599), .A2(new_n613), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n354), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n360), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n366), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n629), .B1(new_n366), .B2(new_n632), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n593), .B(new_n635), .C1(new_n596), .C2(new_n598), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n308), .A2(new_n314), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT95), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n597), .B2(new_n594), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(KEYINPUT100), .A3(new_n593), .A4(new_n635), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n638), .A2(new_n466), .A3(new_n588), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(new_n311), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n633), .A2(new_n634), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n587), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT102), .B(G900), .Z(new_n652));
  AND2_X1   g466(.A1(new_n406), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n404), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n625), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(new_n543), .B(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n400), .A2(new_n544), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n635), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n591), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n656), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n664), .B1(KEYINPUT40), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n310), .A2(new_n306), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n297), .A2(new_n299), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n272), .B2(new_n285), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(G902), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n669), .B1(G472), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n464), .A2(new_n465), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n668), .B(new_n675), .C1(KEYINPUT40), .C2(new_n667), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND4_X1  g491(.A1(new_n464), .A2(new_n465), .A3(new_n609), .A4(new_n656), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n651), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n566), .A2(new_n570), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n575), .B1(new_n682), .B2(new_n577), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n545), .A3(new_n576), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n370), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n617), .B2(new_n618), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NOR2_X1   g503(.A1(new_n625), .A2(new_n613), .ZN(new_n690));
  INV_X1    g504(.A(new_n685), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n311), .A3(new_n369), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND2_X1  g507(.A1(new_n543), .A2(new_n544), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n650), .A3(new_n685), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n674), .A2(new_n311), .A3(new_n695), .A4(new_n409), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(new_n304), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n290), .B2(new_n272), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n295), .B1(new_n699), .B2(new_n300), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n641), .B1(new_n308), .B2(new_n314), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n366), .A2(new_n361), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n684), .A2(new_n610), .A3(new_n545), .A4(new_n576), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n662), .B1(new_n541), .B2(new_n542), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n464), .A3(new_n465), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NOR2_X1   g521(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n679), .A2(new_n695), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT104), .B(G125), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G27));
  NAND3_X1  g525(.A1(new_n311), .A2(new_n366), .A3(new_n361), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT106), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n541), .A2(new_n544), .A3(new_n542), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n591), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n678), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n311), .A2(new_n369), .A3(new_n716), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n679), .A2(new_n721), .A3(KEYINPUT105), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n678), .B2(new_n720), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n714), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n658), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  OAI21_X1  g543(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT107), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n546), .B1(new_n730), .B2(new_n731), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n584), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n576), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT108), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n545), .A3(new_n666), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  INV_X1    g557(.A(new_n465), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT94), .B1(new_n624), .B2(new_n449), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n609), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n674), .A2(KEYINPUT43), .A3(new_n609), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n650), .B1(new_n643), .B2(new_n593), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n715), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(KEYINPUT44), .A3(new_n751), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n742), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  NAND4_X1  g572(.A1(new_n679), .A2(new_n649), .A3(new_n368), .A4(new_n755), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n736), .B1(new_n763), .B2(new_n738), .ZN(new_n764));
  INV_X1    g578(.A(new_n545), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n545), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n759), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n318), .ZN(G42));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n715), .A2(new_n685), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n673), .A2(new_n369), .A3(new_n405), .A4(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n464), .A2(new_n465), .A3(new_n609), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n401), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n404), .B1(new_n748), .B2(new_n749), .ZN(new_n775));
  INV_X1    g589(.A(new_n708), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n702), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n694), .A2(new_n685), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n775), .A2(new_n713), .A3(new_n771), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT48), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT117), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT117), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT48), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n713), .A3(new_n787), .A4(new_n771), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n770), .B(new_n781), .C1(new_n786), .C2(new_n791), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n784), .A2(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n793));
  INV_X1    g607(.A(new_n781), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT118), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n684), .A2(new_n576), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n765), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n766), .A2(new_n767), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n778), .A2(new_n715), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(KEYINPUT51), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n674), .A2(new_n747), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT114), .B1(new_n772), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n775), .A2(new_n771), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n708), .A2(new_n635), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n798), .B2(new_n799), .ZN(new_n810));
  INV_X1    g624(.A(new_n544), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n691), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n661), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n778), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT50), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n802), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n810), .A3(new_n816), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n792), .A2(new_n795), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n696), .A2(new_n706), .A3(new_n692), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n687), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n599), .A2(new_n613), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n400), .B1(new_n744), .B2(new_n745), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n773), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n410), .B(new_n587), .C1(new_n464), .C2(new_n465), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n824), .A2(new_n826), .B1(new_n827), .B2(new_n371), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT109), .B1(new_n828), .B2(new_n645), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n464), .A2(new_n465), .A3(new_n609), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n464), .A2(new_n465), .B1(new_n399), .B2(new_n396), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(KEYINPUT109), .A2(new_n832), .A3(new_n645), .A4(new_n589), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n823), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n400), .A2(new_n657), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n311), .A2(new_n624), .A3(new_n449), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n678), .B2(new_n776), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n717), .A2(new_n650), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n728), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n726), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n659), .A2(new_n709), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n656), .B(KEYINPUT111), .Z(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n848), .B(new_n359), .C1(new_n360), .C2(new_n631), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT112), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(KEYINPUT112), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n665), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n673), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n746), .A3(new_n705), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n845), .A2(new_n846), .A3(new_n680), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n659), .A3(new_n680), .A4(new_n709), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n843), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT110), .B1(new_n834), .B2(new_n842), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n687), .A2(new_n822), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n832), .A2(new_n645), .A3(new_n589), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT109), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n832), .A2(new_n645), .A3(new_n589), .A4(KEYINPUT109), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n840), .B1(new_n725), .B2(new_n719), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n858), .B1(new_n862), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n821), .B(new_n861), .C1(new_n872), .C2(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT113), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n875), .B2(new_n859), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n844), .B2(KEYINPUT52), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n858), .B(new_n877), .C1(new_n862), .C2(new_n871), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n866), .A2(new_n867), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n869), .A2(new_n870), .A3(new_n880), .A4(new_n823), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n859), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n821), .A4(new_n861), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n820), .A2(new_n874), .A3(new_n879), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  INV_X1    g703(.A(new_n796), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT49), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n702), .A2(new_n811), .A3(new_n765), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n890), .A2(KEYINPUT49), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n661), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n674), .A3(new_n609), .A4(new_n673), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n889), .A2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n267), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n861), .ZN(new_n899));
  OAI211_X1 g713(.A(G210), .B(G902), .C1(new_n876), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n504), .A2(new_n508), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n520), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n898), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(KEYINPUT119), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n885), .A2(new_n861), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n909), .A3(G210), .A4(G902), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n906), .A2(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n584), .B(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n821), .B1(new_n885), .B2(new_n861), .ZN(new_n915));
  INV_X1    g729(.A(new_n873), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n683), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n876), .A2(new_n899), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n314), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n733), .A3(new_n734), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n898), .B1(new_n919), .B2(new_n922), .ZN(G54));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n456), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n920), .A2(new_n314), .A3(new_n459), .A4(new_n924), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n898), .ZN(G60));
  NAND3_X1  g742(.A1(new_n874), .A2(new_n879), .A3(new_n887), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n606), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n606), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n915), .B2(new_n916), .ZN(new_n934));
  INV_X1    g748(.A(new_n898), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n932), .A2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT120), .Z(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n348), .B(new_n356), .C1(new_n920), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n885), .B2(new_n861), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n898), .B1(new_n943), .B2(new_n631), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT121), .B1(new_n943), .B2(new_n631), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n942), .B(new_n944), .C1(new_n945), .C2(KEYINPUT61), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n631), .B(new_n940), .C1(new_n876), .C2(new_n899), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n935), .C1(new_n943), .C2(new_n357), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT61), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G66));
  NAND2_X1  g766(.A1(new_n834), .A2(new_n267), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  INV_X1    g768(.A(new_n407), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(G224), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(KEYINPUT122), .B2(new_n953), .ZN(new_n959));
  INV_X1    g773(.A(G898), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n903), .B1(new_n960), .B2(G953), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  AND3_X1   g776(.A1(new_n713), .A2(new_n746), .A3(new_n705), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n742), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n728), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(new_n768), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n844), .B1(new_n651), .B2(new_n679), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n726), .A3(new_n757), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n275), .A2(new_n277), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n452), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(G900), .B2(G953), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n975));
  AOI22_X1  g789(.A1(new_n969), .A2(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n974), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n971), .B(KEYINPUT123), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n666), .B(new_n721), .C1(new_n826), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n981), .B2(new_n826), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n768), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n845), .A2(new_n676), .A3(new_n680), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n967), .A2(new_n987), .A3(new_n676), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n984), .A2(new_n757), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n980), .B1(new_n990), .B2(G953), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n976), .A2(new_n978), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n978), .B1(new_n976), .B2(new_n991), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n968), .B2(new_n834), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n279), .A2(new_n273), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n898), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n876), .A2(new_n878), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n297), .A2(new_n299), .A3(new_n280), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n996), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n996), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n990), .B2(new_n868), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n279), .A2(new_n273), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT127), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n989), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n996), .B1(new_n1009), .B2(new_n834), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n279), .A4(new_n273), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1003), .B1(new_n1007), .B2(new_n1012), .ZN(G57));
endmodule


