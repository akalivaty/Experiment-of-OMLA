

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733;

  OR2_X1 U373 ( .A1(n702), .A2(G902), .ZN(n429) );
  XOR2_X1 U374 ( .A(n433), .B(KEYINPUT89), .Z(n609) );
  NOR2_X1 U375 ( .A1(n541), .A2(n542), .ZN(n637) );
  NAND2_X2 U376 ( .A1(n612), .A2(n611), .ZN(n699) );
  NOR2_X2 U377 ( .A1(n416), .A2(n351), .ZN(n720) );
  XNOR2_X1 U378 ( .A(n417), .B(KEYINPUT48), .ZN(n416) );
  NOR2_X1 U379 ( .A1(n577), .A2(n603), .ZN(n385) );
  NOR2_X1 U380 ( .A1(n577), .A2(n590), .ZN(n386) );
  XNOR2_X1 U381 ( .A(n430), .B(n456), .ZN(n444) );
  XNOR2_X1 U382 ( .A(n503), .B(KEYINPUT4), .ZN(n481) );
  NAND2_X1 U383 ( .A1(n437), .A2(n436), .ZN(n477) );
  XOR2_X1 U384 ( .A(KEYINPUT66), .B(G101), .Z(n462) );
  XNOR2_X1 U385 ( .A(n481), .B(n455), .ZN(n461) );
  INV_X1 U386 ( .A(G134), .ZN(n453) );
  XNOR2_X1 U387 ( .A(n711), .B(n462), .ZN(n480) );
  XNOR2_X1 U388 ( .A(n468), .B(n378), .ZN(n664) );
  INV_X1 U389 ( .A(G472), .ZN(n378) );
  NOR2_X1 U390 ( .A1(n622), .A2(G902), .ZN(n468) );
  OR2_X1 U391 ( .A1(n615), .A2(G902), .ZN(n397) );
  XNOR2_X1 U392 ( .A(n401), .B(n399), .ZN(n517) );
  XNOR2_X1 U393 ( .A(n516), .B(n400), .ZN(n399) );
  OR2_X1 U394 ( .A1(n609), .A2(n607), .ZN(n612) );
  XNOR2_X1 U395 ( .A(n374), .B(n372), .ZN(n696) );
  XNOR2_X1 U396 ( .A(n483), .B(n375), .ZN(n374) );
  INV_X1 U397 ( .A(n710), .ZN(n372) );
  XNOR2_X1 U398 ( .A(n376), .B(n481), .ZN(n375) );
  NOR2_X1 U399 ( .A1(n596), .A2(n648), .ZN(n368) );
  OR2_X1 U400 ( .A1(n577), .A2(n384), .ZN(n578) );
  XOR2_X1 U401 ( .A(G146), .B(KEYINPUT5), .Z(n459) );
  AND2_X1 U402 ( .A1(n588), .A2(n419), .ZN(n418) );
  XOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n485) );
  XNOR2_X1 U404 ( .A(n465), .B(KEYINPUT71), .ZN(n466) );
  XNOR2_X1 U405 ( .A(n480), .B(n479), .ZN(n483) );
  XOR2_X1 U406 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n478) );
  XNOR2_X1 U407 ( .A(n717), .B(n398), .ZN(n615) );
  XNOR2_X1 U408 ( .A(n480), .B(n355), .ZN(n398) );
  INV_X1 U409 ( .A(G953), .ZN(n721) );
  INV_X1 U410 ( .A(KEYINPUT39), .ZN(n422) );
  INV_X1 U411 ( .A(KEYINPUT108), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U413 ( .A(KEYINPUT28), .ZN(n571) );
  NOR2_X1 U414 ( .A1(n589), .A2(n570), .ZN(n377) );
  XNOR2_X1 U415 ( .A(n409), .B(n407), .ZN(n542) );
  XNOR2_X1 U416 ( .A(n408), .B(KEYINPUT103), .ZN(n407) );
  OR2_X1 U417 ( .A1(n698), .A2(G902), .ZN(n409) );
  INV_X1 U418 ( .A(G478), .ZN(n408) );
  XNOR2_X1 U419 ( .A(n411), .B(n410), .ZN(n541) );
  XNOR2_X1 U420 ( .A(n519), .B(G475), .ZN(n410) );
  OR2_X1 U421 ( .A1(n697), .A2(G902), .ZN(n411) );
  XNOR2_X1 U422 ( .A(n498), .B(KEYINPUT0), .ZN(n415) );
  XNOR2_X1 U423 ( .A(n371), .B(n358), .ZN(n370) );
  NAND2_X1 U424 ( .A1(n699), .A2(G472), .ZN(n371) );
  NAND2_X1 U425 ( .A1(n699), .A2(G478), .ZN(n427) );
  NAND2_X1 U426 ( .A1(n699), .A2(G475), .ZN(n383) );
  NAND2_X1 U427 ( .A1(n699), .A2(G469), .ZN(n617) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n515) );
  OR2_X1 U429 ( .A1(G902), .A2(G237), .ZN(n493) );
  INV_X1 U430 ( .A(KEYINPUT44), .ZN(n365) );
  XNOR2_X1 U431 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n438) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n505) );
  XNOR2_X1 U433 ( .A(G107), .B(G134), .ZN(n504) );
  XNOR2_X1 U434 ( .A(G116), .B(G122), .ZN(n502) );
  XNOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT101), .ZN(n400) );
  XNOR2_X1 U436 ( .A(G131), .B(G113), .ZN(n516) );
  XNOR2_X1 U437 ( .A(G122), .B(G143), .ZN(n512) );
  XOR2_X1 U438 ( .A(G140), .B(G104), .Z(n513) );
  XNOR2_X1 U439 ( .A(n402), .B(KEYINPUT11), .ZN(n401) );
  NAND2_X1 U440 ( .A1(n515), .A2(G214), .ZN(n402) );
  XOR2_X1 U441 ( .A(n461), .B(n456), .Z(n717) );
  NOR2_X1 U442 ( .A1(n609), .A2(KEYINPUT2), .ZN(n363) );
  XNOR2_X1 U443 ( .A(n482), .B(KEYINPUT91), .ZN(n376) );
  NOR2_X1 U444 ( .A1(n657), .A2(n658), .ZN(n528) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n622) );
  XNOR2_X1 U446 ( .A(n461), .B(n462), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n463), .B(n487), .ZN(n390) );
  INV_X1 U448 ( .A(n645), .ZN(n605) );
  XNOR2_X1 U449 ( .A(n486), .B(n488), .ZN(n373) );
  INV_X1 U450 ( .A(G122), .ZN(n488) );
  XNOR2_X1 U451 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U452 ( .A(G119), .B(G110), .Z(n430) );
  XOR2_X1 U453 ( .A(G140), .B(KEYINPUT69), .Z(n456) );
  NOR2_X1 U454 ( .A1(n546), .A2(n647), .ZN(n531) );
  INV_X1 U455 ( .A(n664), .ZN(n570) );
  XNOR2_X1 U456 ( .A(n450), .B(n353), .ZN(n428) );
  XNOR2_X1 U457 ( .A(n414), .B(KEYINPUT22), .ZN(n536) );
  INV_X1 U458 ( .A(G104), .ZN(n412) );
  XNOR2_X1 U459 ( .A(n421), .B(n420), .ZN(n733) );
  INV_X1 U460 ( .A(KEYINPUT40), .ZN(n420) );
  AND2_X1 U461 ( .A1(n403), .A2(n599), .ZN(n642) );
  XNOR2_X1 U462 ( .A(n406), .B(n404), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n405), .B(KEYINPUT36), .ZN(n404) );
  INV_X1 U464 ( .A(KEYINPUT80), .ZN(n387) );
  AND2_X1 U465 ( .A1(n584), .A2(n574), .ZN(n388) );
  NAND2_X1 U466 ( .A1(n370), .A2(n381), .ZN(n369) );
  INV_X1 U467 ( .A(KEYINPUT122), .ZN(n423) );
  NAND2_X1 U468 ( .A1(n425), .A2(n381), .ZN(n424) );
  XNOR2_X1 U469 ( .A(n427), .B(n426), .ZN(n425) );
  INV_X1 U470 ( .A(KEYINPUT60), .ZN(n379) );
  NAND2_X1 U471 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U472 ( .A(n383), .B(n359), .ZN(n382) );
  XNOR2_X1 U473 ( .A(n617), .B(n616), .ZN(n618) );
  INV_X1 U474 ( .A(KEYINPUT56), .ZN(n393) );
  NOR2_X1 U475 ( .A1(G953), .A2(n693), .ZN(n695) );
  OR2_X1 U476 ( .A1(n646), .A2(n605), .ZN(n351) );
  XOR2_X1 U477 ( .A(KEYINPUT70), .B(G469), .Z(n352) );
  XOR2_X1 U478 ( .A(n452), .B(n451), .Z(n353) );
  AND2_X1 U479 ( .A1(n679), .A2(n363), .ZN(n354) );
  XOR2_X1 U480 ( .A(n457), .B(G146), .Z(n355) );
  XNOR2_X1 U481 ( .A(n466), .B(n467), .ZN(n487) );
  NOR2_X1 U482 ( .A1(n599), .A2(n661), .ZN(n356) );
  AND2_X1 U483 ( .A1(n508), .A2(G221), .ZN(n357) );
  XNOR2_X1 U484 ( .A(n388), .B(n387), .ZN(n577) );
  XOR2_X1 U485 ( .A(n622), .B(n621), .Z(n358) );
  XNOR2_X1 U486 ( .A(n487), .B(n373), .ZN(n710) );
  XNOR2_X1 U487 ( .A(n697), .B(KEYINPUT59), .ZN(n359) );
  XOR2_X1 U488 ( .A(n696), .B(n431), .Z(n360) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(n623), .Z(n361) );
  NOR2_X1 U490 ( .A1(n733), .A2(n732), .ZN(n586) );
  NOR2_X1 U491 ( .A1(n581), .A2(n649), .ZN(n582) );
  NOR2_X1 U492 ( .A1(n618), .A2(n705), .ZN(n620) );
  INV_X1 U493 ( .A(n705), .ZN(n381) );
  NAND2_X1 U494 ( .A1(n362), .A2(n680), .ZN(n681) );
  NAND2_X1 U495 ( .A1(n679), .A2(KEYINPUT2), .ZN(n362) );
  NOR2_X2 U496 ( .A1(n546), .A2(n521), .ZN(n414) );
  NAND2_X1 U497 ( .A1(n535), .A2(n364), .ZN(n552) );
  NAND2_X1 U498 ( .A1(n366), .A2(n365), .ZN(n364) );
  INV_X1 U499 ( .A(n729), .ZN(n366) );
  XNOR2_X1 U500 ( .A(n448), .B(n357), .ZN(n702) );
  XNOR2_X2 U501 ( .A(n367), .B(n415), .ZN(n546) );
  NAND2_X1 U502 ( .A1(n574), .A2(n497), .ZN(n367) );
  XNOR2_X1 U503 ( .A(n368), .B(n496), .ZN(n574) );
  XNOR2_X1 U504 ( .A(n369), .B(n361), .ZN(G57) );
  XNOR2_X1 U505 ( .A(n377), .B(n571), .ZN(n573) );
  XNOR2_X1 U506 ( .A(n380), .B(n379), .ZN(G60) );
  AND2_X1 U507 ( .A1(n590), .A2(n603), .ZN(n384) );
  XNOR2_X2 U508 ( .A(n391), .B(n533), .ZN(n729) );
  NAND2_X1 U509 ( .A1(n392), .A2(n565), .ZN(n391) );
  XNOR2_X1 U510 ( .A(n531), .B(KEYINPUT34), .ZN(n392) );
  XNOR2_X1 U511 ( .A(n394), .B(n393), .ZN(G51) );
  NAND2_X1 U512 ( .A1(n395), .A2(n381), .ZN(n394) );
  XNOR2_X1 U513 ( .A(n396), .B(n360), .ZN(n395) );
  NAND2_X1 U514 ( .A1(n699), .A2(G210), .ZN(n396) );
  XNOR2_X2 U515 ( .A(n397), .B(n352), .ZN(n572) );
  NAND2_X1 U516 ( .A1(n587), .A2(n418), .ZN(n417) );
  NAND2_X1 U517 ( .A1(n597), .A2(n602), .ZN(n406) );
  XNOR2_X2 U518 ( .A(n413), .B(n412), .ZN(n711) );
  XNOR2_X2 U519 ( .A(G110), .B(G107), .ZN(n413) );
  INV_X1 U520 ( .A(n642), .ZN(n419) );
  NAND2_X1 U521 ( .A1(n604), .A2(n637), .ZN(n421) );
  XNOR2_X1 U522 ( .A(n582), .B(n422), .ZN(n604) );
  XNOR2_X1 U523 ( .A(n424), .B(n423), .ZN(G63) );
  INV_X1 U524 ( .A(n698), .ZN(n426) );
  XNOR2_X2 U525 ( .A(n429), .B(n428), .ZN(n661) );
  XNOR2_X1 U526 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U527 ( .A(n477), .B(n438), .ZN(n511) );
  XNOR2_X2 U528 ( .A(n523), .B(KEYINPUT32), .ZN(n730) );
  XNOR2_X1 U529 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n431) );
  XOR2_X1 U530 ( .A(n614), .B(n613), .Z(n432) );
  XNOR2_X1 U531 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U532 ( .A(KEYINPUT74), .ZN(n527) );
  INV_X1 U533 ( .A(n647), .ZN(n689) );
  INV_X1 U534 ( .A(KEYINPUT81), .ZN(n489) );
  XNOR2_X1 U535 ( .A(n615), .B(n432), .ZN(n616) );
  INV_X1 U536 ( .A(KEYINPUT35), .ZN(n533) );
  NOR2_X1 U537 ( .A1(G952), .A2(n721), .ZN(n705) );
  XNOR2_X1 U538 ( .A(n620), .B(n619), .ZN(G54) );
  XNOR2_X1 U539 ( .A(G902), .B(KEYINPUT15), .ZN(n433) );
  NOR2_X1 U540 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n526) );
  XOR2_X1 U541 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n443) );
  INV_X1 U542 ( .A(G146), .ZN(n434) );
  NAND2_X1 U543 ( .A1(G125), .A2(n434), .ZN(n437) );
  INV_X1 U544 ( .A(G125), .ZN(n435) );
  NAND2_X1 U545 ( .A1(n435), .A2(G146), .ZN(n436) );
  XOR2_X1 U546 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n440) );
  XNOR2_X1 U547 ( .A(G128), .B(G137), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n511), .B(n441), .ZN(n442) );
  XNOR2_X1 U550 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n448) );
  NAND2_X1 U552 ( .A1(n721), .A2(G234), .ZN(n447) );
  XNOR2_X1 U553 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n446) );
  XNOR2_X1 U554 ( .A(n447), .B(n446), .ZN(n508) );
  NAND2_X1 U555 ( .A1(G234), .A2(n609), .ZN(n449) );
  XNOR2_X1 U556 ( .A(KEYINPUT20), .B(n449), .ZN(n499) );
  NAND2_X1 U557 ( .A1(n499), .A2(G217), .ZN(n450) );
  XOR2_X1 U558 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n452) );
  XNOR2_X1 U559 ( .A(KEYINPUT78), .B(KEYINPUT97), .ZN(n451) );
  XNOR2_X2 U560 ( .A(G143), .B(G128), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G131), .B(G137), .ZN(n454) );
  NAND2_X1 U562 ( .A1(G227), .A2(n721), .ZN(n457) );
  XNOR2_X2 U563 ( .A(n572), .B(KEYINPUT1), .ZN(n657) );
  NOR2_X1 U564 ( .A1(n661), .A2(n657), .ZN(n469) );
  NAND2_X1 U565 ( .A1(G210), .A2(n515), .ZN(n458) );
  XNOR2_X1 U566 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U567 ( .A(n460), .B(KEYINPUT75), .Z(n463) );
  XNOR2_X1 U568 ( .A(G113), .B(G119), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n464), .B(KEYINPUT3), .ZN(n467) );
  XNOR2_X1 U570 ( .A(G116), .B(KEYINPUT90), .ZN(n465) );
  XOR2_X1 U571 ( .A(KEYINPUT6), .B(n664), .Z(n592) );
  INV_X1 U572 ( .A(n592), .ZN(n537) );
  NAND2_X1 U573 ( .A1(n469), .A2(n537), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n470), .B(KEYINPUT79), .ZN(n522) );
  NOR2_X1 U575 ( .A1(G898), .A2(n721), .ZN(n714) );
  NAND2_X1 U576 ( .A1(G237), .A2(G234), .ZN(n471) );
  XNOR2_X1 U577 ( .A(n471), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U578 ( .A1(G902), .A2(n473), .ZN(n554) );
  INV_X1 U579 ( .A(n554), .ZN(n472) );
  NAND2_X1 U580 ( .A1(n714), .A2(n472), .ZN(n476) );
  NAND2_X1 U581 ( .A1(G952), .A2(n473), .ZN(n474) );
  XOR2_X1 U582 ( .A(KEYINPUT93), .B(n474), .Z(n676) );
  NOR2_X1 U583 ( .A1(G953), .A2(n676), .ZN(n558) );
  INV_X1 U584 ( .A(n558), .ZN(n475) );
  NAND2_X1 U585 ( .A1(n476), .A2(n475), .ZN(n497) );
  NAND2_X1 U586 ( .A1(G224), .A2(n721), .ZN(n482) );
  INV_X1 U587 ( .A(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U588 ( .A1(n696), .A2(n609), .ZN(n492) );
  NAND2_X1 U589 ( .A1(n493), .A2(G210), .ZN(n490) );
  XNOR2_X2 U590 ( .A(n492), .B(n491), .ZN(n596) );
  NAND2_X1 U591 ( .A1(n493), .A2(G214), .ZN(n494) );
  XOR2_X1 U592 ( .A(n494), .B(KEYINPUT92), .Z(n648) );
  XNOR2_X1 U593 ( .A(KEYINPUT19), .B(KEYINPUT64), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n495), .B(KEYINPUT77), .ZN(n496) );
  XNOR2_X1 U595 ( .A(KEYINPUT65), .B(KEYINPUT87), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n501) );
  NAND2_X1 U597 ( .A1(n499), .A2(G221), .ZN(n500) );
  XNOR2_X1 U598 ( .A(n501), .B(n500), .ZN(n660) );
  XOR2_X1 U599 ( .A(n503), .B(n502), .Z(n507) );
  XNOR2_X1 U600 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U601 ( .A(n507), .B(n506), .Z(n510) );
  NAND2_X1 U602 ( .A1(G217), .A2(n508), .ZN(n509) );
  XOR2_X1 U603 ( .A(n510), .B(n509), .Z(n698) );
  XNOR2_X1 U604 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n519) );
  BUF_X1 U605 ( .A(n511), .Z(n718) );
  XNOR2_X1 U606 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U607 ( .A(n718), .B(n514), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n518), .B(n517), .ZN(n697) );
  INV_X1 U609 ( .A(n541), .ZN(n520) );
  NOR2_X1 U610 ( .A1(n542), .A2(n520), .ZN(n650) );
  NAND2_X1 U611 ( .A1(n660), .A2(n650), .ZN(n521) );
  NAND2_X1 U612 ( .A1(n522), .A2(n536), .ZN(n523) );
  INV_X1 U613 ( .A(n657), .ZN(n599) );
  AND2_X1 U614 ( .A1(n536), .A2(n356), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n524), .A2(n570), .ZN(n633) );
  NAND2_X1 U616 ( .A1(n730), .A2(n633), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n526), .B(n525), .ZN(n534) );
  NAND2_X1 U618 ( .A1(n660), .A2(n661), .ZN(n658) );
  XNOR2_X1 U619 ( .A(n528), .B(n527), .ZN(n545) );
  NOR2_X1 U620 ( .A1(n545), .A2(n537), .ZN(n530) );
  XNOR2_X1 U621 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n529) );
  XNOR2_X1 U622 ( .A(n530), .B(n529), .ZN(n647) );
  INV_X1 U623 ( .A(n542), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n541), .A2(n532), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n534), .A2(n729), .ZN(n535) );
  AND2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U627 ( .A(n538), .B(KEYINPUT84), .ZN(n539) );
  AND2_X1 U628 ( .A1(n539), .A2(n657), .ZN(n540) );
  AND2_X1 U629 ( .A1(n661), .A2(n540), .ZN(n624) );
  INV_X1 U630 ( .A(n637), .ZN(n590) );
  NAND2_X1 U631 ( .A1(n542), .A2(n541), .ZN(n603) );
  NAND2_X1 U632 ( .A1(n590), .A2(n603), .ZN(n652) );
  NOR2_X1 U633 ( .A1(n572), .A2(n658), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n563), .A2(n570), .ZN(n543) );
  NOR2_X1 U635 ( .A1(n546), .A2(n543), .ZN(n630) );
  XOR2_X1 U636 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n544) );
  XNOR2_X1 U637 ( .A(KEYINPUT31), .B(n544), .ZN(n548) );
  OR2_X1 U638 ( .A1(n570), .A2(n545), .ZN(n667) );
  NOR2_X1 U639 ( .A1(n546), .A2(n667), .ZN(n547) );
  XOR2_X1 U640 ( .A(n548), .B(n547), .Z(n640) );
  NOR2_X1 U641 ( .A1(n630), .A2(n640), .ZN(n549) );
  NOR2_X1 U642 ( .A1(n384), .A2(n549), .ZN(n550) );
  NOR2_X1 U643 ( .A1(n624), .A2(n550), .ZN(n551) );
  NAND2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X2 U645 ( .A(n553), .B(KEYINPUT45), .ZN(n679) );
  NOR2_X1 U646 ( .A1(G900), .A2(n554), .ZN(n555) );
  NAND2_X1 U647 ( .A1(G953), .A2(n555), .ZN(n556) );
  XOR2_X1 U648 ( .A(KEYINPUT104), .B(n556), .Z(n557) );
  NOR2_X1 U649 ( .A1(n558), .A2(n557), .ZN(n568) );
  XOR2_X1 U650 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n560) );
  INV_X1 U651 ( .A(n648), .ZN(n594) );
  NAND2_X1 U652 ( .A1(n664), .A2(n594), .ZN(n559) );
  XNOR2_X1 U653 ( .A(n560), .B(n559), .ZN(n561) );
  NOR2_X1 U654 ( .A1(n568), .A2(n561), .ZN(n562) );
  NAND2_X1 U655 ( .A1(n563), .A2(n562), .ZN(n581) );
  NOR2_X1 U656 ( .A1(n596), .A2(n581), .ZN(n564) );
  NAND2_X1 U657 ( .A1(n565), .A2(n564), .ZN(n635) );
  NAND2_X1 U658 ( .A1(n384), .A2(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n635), .A2(n566), .ZN(n567) );
  XOR2_X1 U660 ( .A(KEYINPUT82), .B(n567), .Z(n576) );
  NOR2_X1 U661 ( .A1(n661), .A2(n568), .ZN(n569) );
  NAND2_X1 U662 ( .A1(n660), .A2(n569), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n573), .A2(n572), .ZN(n584) );
  NAND2_X1 U664 ( .A1(KEYINPUT47), .A2(n577), .ZN(n575) );
  NAND2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n580) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(n578), .ZN(n579) );
  NOR2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n588) );
  XOR2_X1 U668 ( .A(n596), .B(KEYINPUT38), .Z(n649) );
  NOR2_X1 U669 ( .A1(n648), .A2(n649), .ZN(n653) );
  NAND2_X1 U670 ( .A1(n653), .A2(n650), .ZN(n583) );
  XNOR2_X1 U671 ( .A(n583), .B(KEYINPUT41), .ZN(n688) );
  AND2_X1 U672 ( .A1(n584), .A2(n688), .ZN(n585) );
  XNOR2_X1 U673 ( .A(n585), .B(KEYINPUT42), .ZN(n732) );
  XNOR2_X1 U674 ( .A(n586), .B(KEYINPUT46), .ZN(n587) );
  NOR2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U677 ( .A(KEYINPUT105), .B(n593), .ZN(n595) );
  AND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U679 ( .A(n596), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT106), .B(n597), .Z(n598) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT43), .ZN(n601) );
  NOR2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n646) );
  INV_X1 U684 ( .A(n603), .ZN(n639) );
  NAND2_X1 U685 ( .A1(n639), .A2(n604), .ZN(n645) );
  NAND2_X1 U686 ( .A1(n679), .A2(n720), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  INV_X1 U688 ( .A(n720), .ZN(n677) );
  INV_X1 U689 ( .A(KEYINPUT76), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n677), .B(n608), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n610), .A2(n354), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n614) );
  XNOR2_X1 U693 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n613) );
  INV_X1 U694 ( .A(KEYINPUT121), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n621) );
  XOR2_X1 U696 ( .A(KEYINPUT63), .B(KEYINPUT110), .Z(n623) );
  XOR2_X1 U697 ( .A(G101), .B(n624), .Z(G3) );
  XOR2_X1 U698 ( .A(G104), .B(KEYINPUT111), .Z(n626) );
  NAND2_X1 U699 ( .A1(n630), .A2(n637), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n628) );
  XNOR2_X1 U702 ( .A(G107), .B(KEYINPUT112), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n629) );
  XOR2_X1 U704 ( .A(KEYINPUT26), .B(n629), .Z(n632) );
  NAND2_X1 U705 ( .A1(n630), .A2(n639), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(G9) );
  XNOR2_X1 U707 ( .A(G110), .B(n633), .ZN(G12) );
  XNOR2_X1 U708 ( .A(G128), .B(n385), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT29), .ZN(G30) );
  XNOR2_X1 U710 ( .A(G143), .B(n635), .ZN(G45) );
  XOR2_X1 U711 ( .A(G146), .B(n386), .Z(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT114), .B(n636), .ZN(G48) );
  NAND2_X1 U713 ( .A1(n640), .A2(n637), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n638), .B(G113), .ZN(G15) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(G116), .ZN(G18) );
  XOR2_X1 U717 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U718 ( .A(G125), .B(n642), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G27) );
  XNOR2_X1 U720 ( .A(G134), .B(n645), .ZN(G36) );
  XOR2_X1 U721 ( .A(G140), .B(n646), .Z(G42) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n689), .A2(n656), .ZN(n672) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT51), .B(n669), .Z(n670) );
  NAND2_X1 U735 ( .A1(n688), .A2(n670), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U737 ( .A(n673), .B(KEYINPUT52), .ZN(n674) );
  XOR2_X1 U738 ( .A(KEYINPUT116), .B(n674), .Z(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n687) );
  INV_X1 U740 ( .A(KEYINPUT83), .ZN(n680) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(n680), .Z(n678) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n681), .A2(n720), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n679), .A2(KEYINPUT2), .ZN(n684) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n692) );
  AND2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(KEYINPUT117), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U751 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n695), .B(n694), .ZN(G75) );
  XOR2_X1 U753 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n701) );
  NAND2_X1 U754 ( .A1(n699), .A2(G217), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n705), .A2(n704), .ZN(G66) );
  NAND2_X1 U758 ( .A1(n721), .A2(n679), .ZN(n709) );
  NAND2_X1 U759 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U760 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U761 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n716) );
  XNOR2_X1 U763 ( .A(n710), .B(G101), .ZN(n712) );
  XNOR2_X1 U764 ( .A(n711), .B(n712), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(n715), .ZN(G69) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U768 ( .A(n719), .B(KEYINPUT125), .Z(n724) );
  XOR2_X1 U769 ( .A(n724), .B(n720), .Z(n722) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT126), .ZN(n728) );
  XNOR2_X1 U772 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(n726), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G122), .B(n729), .ZN(G24) );
  XOR2_X1 U777 ( .A(n730), .B(G119), .Z(n731) );
  XNOR2_X1 U778 ( .A(KEYINPUT127), .B(n731), .ZN(G21) );
  XOR2_X1 U779 ( .A(G137), .B(n732), .Z(G39) );
  XOR2_X1 U780 ( .A(n733), .B(G131), .Z(G33) );
endmodule

