

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n542), .A2(G2104), .ZN(n881) );
  AND2_X1 U550 ( .A1(n741), .A2(n969), .ZN(n515) );
  INV_X1 U551 ( .A(KEYINPUT96), .ZN(n681) );
  XNOR2_X1 U552 ( .A(n723), .B(n681), .ZN(n707) );
  INV_X1 U553 ( .A(KEYINPUT31), .ZN(n719) );
  INV_X1 U554 ( .A(n980), .ZN(n748) );
  INV_X1 U555 ( .A(KEYINPUT103), .ZN(n759) );
  OR2_X1 U556 ( .A1(n676), .A2(n675), .ZN(n773) );
  NOR2_X1 U557 ( .A1(n677), .A2(G1384), .ZN(n774) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n538) );
  NAND2_X1 U559 ( .A1(n882), .A2(G138), .ZN(n540) );
  NOR2_X1 U560 ( .A1(G2104), .A2(n542), .ZN(n878) );
  NOR2_X1 U561 ( .A1(G651), .A2(n608), .ZN(n643) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n521), .Z(n644) );
  NOR2_X1 U563 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U564 ( .A1(n639), .A2(G89), .ZN(n516) );
  XNOR2_X1 U565 ( .A(n516), .B(KEYINPUT4), .ZN(n518) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n608) );
  INV_X1 U567 ( .A(G651), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n608), .A2(n520), .ZN(n638) );
  NAND2_X1 U569 ( .A1(G76), .A2(n638), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n519), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U572 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G51), .A2(n643), .ZN(n523) );
  NOR2_X1 U574 ( .A1(G543), .A2(n520), .ZN(n521) );
  NAND2_X1 U575 ( .A1(G63), .A2(n644), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U577 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U579 ( .A(KEYINPUT7), .B(n528), .ZN(G168) );
  XOR2_X1 U580 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U581 ( .A(KEYINPUT9), .B(KEYINPUT67), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G77), .A2(n638), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G90), .A2(n639), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n532), .B(n531), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n644), .A2(G64), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n533), .B(KEYINPUT66), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G52), .A2(n643), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(G171) );
  INV_X1 U591 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G102), .A2(n881), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XNOR2_X2 U594 ( .A(n539), .B(n538), .ZN(n882) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n546) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U597 ( .A1(G114), .A2(n877), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G126), .A2(n878), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n677) );
  BUF_X1 U601 ( .A(n677), .Z(G164) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G120), .ZN(G236) );
  INV_X1 U605 ( .A(G69), .ZN(G235) );
  INV_X1 U606 ( .A(G108), .ZN(G238) );
  NAND2_X1 U607 ( .A1(G91), .A2(n639), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G65), .A2(n644), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G53), .A2(n643), .ZN(n549) );
  XNOR2_X1 U611 ( .A(KEYINPUT69), .B(n549), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n638), .A2(G78), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U615 ( .A1(n882), .A2(G137), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G101), .A2(n881), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT23), .B(n554), .Z(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n675) );
  NAND2_X1 U619 ( .A1(G125), .A2(n878), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G113), .A2(n877), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n673) );
  NOR2_X1 U622 ( .A1(n675), .A2(n673), .ZN(G160) );
  NAND2_X1 U623 ( .A1(G94), .A2(G452), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(n559), .Z(G173) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT70), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT10), .B(n561), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n815) );
  NAND2_X1 U629 ( .A1(n815), .A2(G567), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT71), .ZN(n563) );
  XNOR2_X1 U631 ( .A(KEYINPUT11), .B(n563), .ZN(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n644), .ZN(n564) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n564), .Z(n571) );
  NAND2_X1 U634 ( .A1(G81), .A2(n639), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n565), .B(KEYINPUT72), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G68), .A2(n638), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(n569), .Z(n570) );
  NOR2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n643), .A2(G43), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n966) );
  INV_X1 U643 ( .A(G860), .ZN(n588) );
  OR2_X1 U644 ( .A1(n966), .A2(n588), .ZN(G153) );
  XNOR2_X1 U645 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n574) );
  XOR2_X1 U647 ( .A(KEYINPUT74), .B(n574), .Z(n584) );
  NAND2_X1 U648 ( .A1(G54), .A2(n643), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G79), .A2(n638), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G92), .A2(n639), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G66), .A2(n644), .ZN(n577) );
  XNOR2_X1 U653 ( .A(KEYINPUT75), .B(n577), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X2 U656 ( .A(n582), .B(KEYINPUT15), .ZN(n973) );
  NOR2_X1 U657 ( .A1(n973), .A2(G868), .ZN(n583) );
  NOR2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U659 ( .A(KEYINPUT76), .B(n585), .Z(G284) );
  INV_X1 U660 ( .A(G868), .ZN(n656) );
  NOR2_X1 U661 ( .A1(G286), .A2(n656), .ZN(n587) );
  NOR2_X1 U662 ( .A1(G868), .A2(G299), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n587), .A2(n586), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n588), .A2(G559), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n589), .A2(n973), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT16), .ZN(n591) );
  XNOR2_X1 U667 ( .A(KEYINPUT78), .B(n591), .ZN(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n966), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G868), .A2(n973), .ZN(n592) );
  NOR2_X1 U670 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G99), .A2(n881), .ZN(n596) );
  NAND2_X1 U673 ( .A1(G111), .A2(n877), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT79), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G135), .A2(n882), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n878), .A2(G123), .ZN(n600) );
  XOR2_X1 U679 ( .A(KEYINPUT18), .B(n600), .Z(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n917) );
  XNOR2_X1 U681 ( .A(n917), .B(G2096), .ZN(n604) );
  INV_X1 U682 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G49), .A2(n643), .ZN(n606) );
  NAND2_X1 U685 ( .A1(G74), .A2(G651), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n644), .A2(n607), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n608), .A2(G87), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G288) );
  NAND2_X1 U690 ( .A1(G73), .A2(n638), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT2), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G48), .A2(n643), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G61), .A2(n644), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G86), .A2(n639), .ZN(n614) );
  XNOR2_X1 U696 ( .A(KEYINPUT85), .B(n614), .ZN(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT86), .B(n619), .ZN(G305) );
  NAND2_X1 U700 ( .A1(G50), .A2(n643), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G62), .A2(n644), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT87), .B(n622), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G75), .A2(n638), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G88), .A2(n639), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U707 ( .A(KEYINPUT88), .B(n625), .Z(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(G303) );
  INV_X1 U709 ( .A(G303), .ZN(G166) );
  NAND2_X1 U710 ( .A1(G72), .A2(n638), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G85), .A2(n639), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G60), .A2(n644), .ZN(n630) );
  XNOR2_X1 U714 ( .A(KEYINPUT65), .B(n630), .ZN(n631) );
  NOR2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n643), .A2(G47), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(G290) );
  XNOR2_X1 U718 ( .A(n966), .B(KEYINPUT80), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n973), .A2(G559), .ZN(n635) );
  XNOR2_X1 U720 ( .A(n636), .B(n635), .ZN(n819) );
  XOR2_X1 U721 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n637) );
  XNOR2_X1 U722 ( .A(G288), .B(n637), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G80), .A2(n638), .ZN(n641) );
  NAND2_X1 U724 ( .A1(G93), .A2(n639), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U726 ( .A(KEYINPUT82), .B(n642), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G55), .A2(n643), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G67), .A2(n644), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U731 ( .A(KEYINPUT83), .B(n649), .ZN(n822) );
  XNOR2_X1 U732 ( .A(n650), .B(n822), .ZN(n652) );
  XNOR2_X1 U733 ( .A(G305), .B(G166), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U735 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(G299), .ZN(n845) );
  XNOR2_X1 U737 ( .A(n819), .B(n845), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n655), .A2(G868), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n656), .A2(n822), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G235), .A2(G236), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(KEYINPUT91), .ZN(n664) );
  NOR2_X1 U749 ( .A1(G238), .A2(n664), .ZN(n665) );
  NAND2_X1 U750 ( .A1(G57), .A2(n665), .ZN(n825) );
  NAND2_X1 U751 ( .A1(n825), .A2(G567), .ZN(n671) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U754 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U755 ( .A1(G96), .A2(n668), .ZN(n824) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n824), .ZN(n669) );
  XNOR2_X1 U757 ( .A(KEYINPUT90), .B(n669), .ZN(n670) );
  NAND2_X1 U758 ( .A1(n671), .A2(n670), .ZN(n826) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U760 ( .A1(n826), .A2(n672), .ZN(n818) );
  NAND2_X1 U761 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(n673), .ZN(n674) );
  NAND2_X1 U763 ( .A1(G40), .A2(n674), .ZN(n676) );
  INV_X1 U764 ( .A(n773), .ZN(n678) );
  NAND2_X2 U765 ( .A1(n678), .A2(n774), .ZN(n723) );
  NAND2_X1 U766 ( .A1(G8), .A2(n723), .ZN(n755) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n679) );
  XOR2_X1 U768 ( .A(n679), .B(KEYINPUT24), .Z(n680) );
  NOR2_X1 U769 ( .A1(n755), .A2(n680), .ZN(n762) );
  NAND2_X1 U770 ( .A1(n707), .A2(G2067), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G1348), .A2(n723), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n683), .A2(n682), .ZN(n690) );
  INV_X1 U773 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U774 ( .A1(n723), .A2(n942), .ZN(n685) );
  XOR2_X1 U775 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n684) );
  XNOR2_X1 U776 ( .A(n685), .B(n684), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n723), .A2(G1341), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U779 ( .A1(n966), .A2(n688), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n973), .A2(n692), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT97), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n973), .A2(n692), .ZN(n693) );
  NOR2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n707), .A2(G2072), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT27), .B(n695), .Z(n698) );
  INV_X1 U787 ( .A(n707), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n696), .A2(G1956), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U790 ( .A1(G299), .A2(n702), .ZN(n699) );
  XNOR2_X1 U791 ( .A(n699), .B(KEYINPUT98), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U793 ( .A1(G299), .A2(n702), .ZN(n703) );
  XOR2_X1 U794 ( .A(KEYINPUT28), .B(n703), .Z(n704) );
  NOR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U796 ( .A(n706), .B(KEYINPUT29), .ZN(n711) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NAND2_X1 U798 ( .A1(n707), .A2(n941), .ZN(n709) );
  INV_X1 U799 ( .A(G1961), .ZN(n990) );
  NAND2_X1 U800 ( .A1(n990), .A2(n723), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n716) );
  NAND2_X1 U802 ( .A1(G171), .A2(n716), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n722) );
  NOR2_X1 U804 ( .A1(G1966), .A2(n755), .ZN(n733) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n723), .ZN(n732) );
  NOR2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n712) );
  NAND2_X1 U807 ( .A1(G8), .A2(n712), .ZN(n713) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n713), .ZN(n714) );
  NOR2_X1 U809 ( .A1(G168), .A2(n714), .ZN(n715) );
  XOR2_X1 U810 ( .A(KEYINPUT99), .B(n715), .Z(n718) );
  NOR2_X1 U811 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n736) );
  NAND2_X1 U815 ( .A1(n736), .A2(G286), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n723), .ZN(n724) );
  XNOR2_X1 U817 ( .A(KEYINPUT101), .B(n724), .ZN(n727) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n755), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G166), .A2(n725), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT32), .ZN(n739) );
  AND2_X1 U824 ( .A1(G8), .A2(n732), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U827 ( .A(KEYINPUT100), .B(n737), .Z(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n752) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n745) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n745), .A2(n740), .ZN(n970) );
  NAND2_X1 U832 ( .A1(n752), .A2(n970), .ZN(n742) );
  INV_X1 U833 ( .A(n755), .ZN(n741) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NAND2_X1 U835 ( .A1(n742), .A2(n515), .ZN(n744) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n743) );
  NAND2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n750) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n980) );
  NAND2_X1 U839 ( .A1(n745), .A2(KEYINPUT33), .ZN(n746) );
  NOR2_X1 U840 ( .A1(n755), .A2(n746), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT102), .ZN(n758) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U845 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n752), .A2(n754), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(n759), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n795) );
  XNOR2_X1 U851 ( .A(KEYINPUT37), .B(G2067), .ZN(n808) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G104), .A2(n881), .ZN(n764) );
  NAND2_X1 U854 ( .A1(G140), .A2(n882), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U856 ( .A(n766), .B(n765), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G116), .A2(n877), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G128), .A2(n878), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U860 ( .A(KEYINPUT35), .B(n769), .Z(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U862 ( .A(KEYINPUT36), .B(n772), .ZN(n872) );
  NOR2_X1 U863 ( .A1(n808), .A2(n872), .ZN(n921) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n810) );
  NAND2_X1 U865 ( .A1(n921), .A2(n810), .ZN(n775) );
  XOR2_X1 U866 ( .A(KEYINPUT93), .B(n775), .Z(n805) );
  NAND2_X1 U867 ( .A1(G95), .A2(n881), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G131), .A2(n882), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G107), .A2(n877), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G119), .A2(n878), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n862) );
  INV_X1 U874 ( .A(G1991), .ZN(n945) );
  NOR2_X1 U875 ( .A1(n862), .A2(n945), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G117), .A2(n877), .ZN(n783) );
  NAND2_X1 U877 ( .A1(G129), .A2(n878), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U879 ( .A(KEYINPUT94), .B(n784), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n881), .A2(G105), .ZN(n785) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n882), .A2(G141), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n888) );
  AND2_X1 U885 ( .A1(n888), .A2(G1996), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n923) );
  INV_X1 U887 ( .A(n810), .ZN(n792) );
  NOR2_X1 U888 ( .A1(n923), .A2(n792), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT95), .B(n800), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n805), .A2(n793), .ZN(n794) );
  NOR2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n797) );
  XNOR2_X1 U892 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U893 ( .A1(n977), .A2(n810), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n813) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n888), .ZN(n929) );
  AND2_X1 U896 ( .A1(n945), .A2(n862), .ZN(n918) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U898 ( .A1(n918), .A2(n798), .ZN(n799) );
  NOR2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U900 ( .A(n801), .B(KEYINPUT104), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n929), .A2(n802), .ZN(n803) );
  XOR2_X1 U902 ( .A(n803), .B(KEYINPUT39), .Z(n804) );
  XNOR2_X1 U903 ( .A(KEYINPUT105), .B(n804), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U905 ( .A(n807), .B(KEYINPUT106), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n808), .A2(n872), .ZN(n933) );
  NAND2_X1 U907 ( .A1(n809), .A2(n933), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U913 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(G188) );
  XNOR2_X1 U917 ( .A(KEYINPUT81), .B(KEYINPUT84), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n819), .A2(G860), .ZN(n820) );
  XNOR2_X1 U919 ( .A(n821), .B(n820), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(G145) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  NOR2_X1 U922 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n826), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2100), .B(G2096), .Z(n828) );
  XNOR2_X1 U926 ( .A(KEYINPUT42), .B(G2678), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2090), .Z(n830) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U931 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2084), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1956), .B(G1961), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1981), .B(G1966), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(G1976), .B(G1971), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(KEYINPUT109), .B(G2474), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U943 ( .A(G1986), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G229) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT115), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n966), .B(G286), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n973), .B(G171), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  NOR2_X1 U950 ( .A1(G37), .A2(n850), .ZN(G397) );
  NAND2_X1 U951 ( .A1(G100), .A2(n881), .ZN(n852) );
  NAND2_X1 U952 ( .A1(G112), .A2(n877), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n858) );
  NAND2_X1 U954 ( .A1(G124), .A2(n878), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G136), .A2(n882), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n854), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U959 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n860) );
  XNOR2_X1 U961 ( .A(G162), .B(KEYINPUT113), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n876) );
  NAND2_X1 U964 ( .A1(G103), .A2(n881), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G139), .A2(n882), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n878), .A2(G127), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n877), .A2(G115), .ZN(n865) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n865), .Z(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U972 ( .A(n869), .B(n868), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n912) );
  XNOR2_X1 U974 ( .A(n872), .B(n912), .ZN(n874) );
  XNOR2_X1 U975 ( .A(G164), .B(G160), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n892) );
  NAND2_X1 U978 ( .A1(G118), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U987 ( .A(n917), .B(n890), .Z(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U989 ( .A1(G37), .A2(n893), .ZN(n894) );
  XNOR2_X1 U990 ( .A(KEYINPUT114), .B(n894), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G2451), .B(G2427), .ZN(n904) );
  XOR2_X1 U992 ( .A(G2430), .B(G2443), .Z(n896) );
  XNOR2_X1 U993 ( .A(G2435), .B(KEYINPUT107), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U995 ( .A(G2438), .B(G2454), .Z(n898) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U999 ( .A(G2446), .B(KEYINPUT108), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(n905), .A2(G14), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G57), .ZN(G237) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n938) );
  XNOR2_X1 U1013 ( .A(G164), .B(G2078), .ZN(n915) );
  XOR2_X1 U1014 ( .A(G2072), .B(n912), .Z(n913) );
  XNOR2_X1 U1015 ( .A(KEYINPUT119), .B(n913), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT50), .ZN(n936) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(KEYINPUT117), .B(n919), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT118), .B(n927), .Z(n932) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT51), .B(n930), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n938), .B(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n939), .B(KEYINPUT52), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(G29), .ZN(n1019) );
  XOR2_X1 U1035 ( .A(n941), .B(G27), .Z(n944) );
  XOR2_X1 U1036 ( .A(n942), .B(G32), .Z(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n955) );
  XNOR2_X1 U1038 ( .A(n945), .B(G25), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT122), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G2072), .B(KEYINPUT123), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G33), .B(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT124), .B(n951), .Z(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(KEYINPUT53), .ZN(n959) );
  XOR2_X1 U1049 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n957), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1054 ( .A(KEYINPUT125), .B(n962), .Z(n963) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n963), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n964), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n965), .A2(G11), .ZN(n1017) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XOR2_X1 U1059 ( .A(G171), .B(G1961), .Z(n968) );
  XNOR2_X1 U1060 ( .A(n966), .B(G1341), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n987) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(G1956), .B(G299), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n979) );
  XNOR2_X1 U1065 ( .A(n973), .B(G1348), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n985) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n982), .B(KEYINPUT126), .ZN(n983) );
  XOR2_X1 U1073 ( .A(KEYINPUT57), .B(n983), .Z(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n1015) );
  INV_X1 U1077 ( .A(G16), .ZN(n1013) );
  XNOR2_X1 U1078 ( .A(G5), .B(n990), .ZN(n1003) );
  XOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .Z(n991) );
  XNOR2_X1 U1080 ( .A(G4), .B(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G20), .B(G1956), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G19), .B(G1341), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT127), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT60), .B(n999), .Z(n1001) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G21), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

