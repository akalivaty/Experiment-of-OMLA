//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT64), .Z(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G238), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n217), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT68), .B(G45), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT76), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT13), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n248), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  MUX2_X1   g0061(.A(new_n261), .B(new_n233), .S(G1698), .Z(new_n262));
  NAND2_X1  g0062(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n260), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n256), .A2(new_n213), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n259), .A2(G238), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n253), .A2(new_n254), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n254), .B1(new_n253), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g0072(.A(G169), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n274));
  INV_X1    g0074(.A(new_n272), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G169), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n270), .A2(KEYINPUT77), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT77), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n253), .A2(new_n269), .A3(new_n280), .A4(new_n254), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n279), .A2(new_n275), .A3(G179), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n274), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n213), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n213), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n207), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G20), .A3(new_n291), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n206), .A2(G20), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT71), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n285), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n298), .B(new_n302), .C1(new_n291), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n283), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n276), .B2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n279), .A2(new_n275), .A3(new_n281), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n257), .A2(new_n258), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n252), .B1(new_n317), .B2(new_n261), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G222), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT69), .B(G223), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT3), .B(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n293), .B2(new_n323), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n318), .B1(new_n325), .B2(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n313), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G200), .B2(new_n326), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT10), .B1(new_n328), .B2(KEYINPUT75), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n294), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n289), .B1(new_n202), .B2(new_n307), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n289), .A2(new_n307), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G50), .A3(new_n305), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT9), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n337), .A2(new_n328), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n329), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n218), .A2(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n319), .A2(G232), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n266), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(G107), .B2(new_n266), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n257), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G244), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n252), .B1(new_n317), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(G179), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(G169), .B1(new_n344), .B2(new_n347), .ZN(new_n350));
  INV_X1    g0150(.A(new_n331), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n353), .A2(KEYINPUT73), .A3(new_n294), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT73), .B1(new_n353), .B2(new_n294), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n285), .ZN(new_n357));
  MUX2_X1   g0157(.A(new_n306), .B(new_n309), .S(G77), .Z(new_n358));
  AOI22_X1  g0158(.A1(new_n349), .A2(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n345), .A2(new_n313), .A3(new_n348), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n344), .B2(new_n347), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n360), .A2(new_n366), .A3(KEYINPUT74), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n359), .B2(new_n365), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n326), .A2(G179), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n326), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n336), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n367), .A2(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n316), .A2(new_n339), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n304), .A2(new_n331), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n334), .A2(new_n379), .B1(new_n307), .B2(new_n331), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n264), .A2(KEYINPUT79), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT80), .A4(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n263), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT80), .B1(new_n387), .B2(G33), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n207), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT7), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n207), .C1(new_n386), .C2(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(G68), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n291), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n201), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n290), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n266), .B2(new_n207), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n265), .B1(new_n387), .B2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n391), .A2(G20), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n399), .B1(new_n404), .B2(new_n291), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n406), .B1(new_n213), .B2(new_n284), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n381), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n382), .A2(new_n384), .A3(G33), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT80), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n319), .A2(G223), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n261), .B2(new_n319), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n411), .A2(new_n263), .A3(new_n385), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n257), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n252), .B1(new_n317), .B2(new_n233), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n363), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(G190), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT17), .B1(new_n408), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n371), .B1(new_n416), .B2(new_n417), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n419), .B2(G179), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT18), .B1(new_n408), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n416), .A2(G179), .A3(new_n417), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n371), .B2(new_n419), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n391), .B1(new_n323), .B2(G20), .ZN(new_n430));
  INV_X1    g0230(.A(new_n265), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n382), .A2(new_n384), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n255), .ZN(new_n433));
  INV_X1    g0233(.A(new_n403), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n398), .B1(new_n435), .B2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n285), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n291), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n398), .B1(new_n438), .B2(new_n392), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n439), .B2(KEYINPUT16), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n427), .B(new_n429), .C1(new_n440), .C2(new_n381), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n426), .A2(new_n441), .A3(KEYINPUT81), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT81), .B1(new_n426), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n423), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n206), .B(G45), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT84), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n450));
  OAI211_X1 g0250(.A(G274), .B(new_n450), .C1(new_n256), .C2(new_n213), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n450), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n445), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n268), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n449), .A2(new_n452), .B1(new_n455), .B2(G257), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n457), .A2(new_n346), .A3(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(G250), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n319), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n323), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n346), .A2(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n411), .A2(new_n263), .A3(new_n385), .A4(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(new_n457), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n456), .B1(new_n466), .B2(new_n257), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n363), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G190), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT6), .A2(G97), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n470), .A2(new_n473), .A3(G107), .ZN(new_n474));
  XOR2_X1   g0274(.A(G97), .B(G107), .Z(new_n475));
  OAI22_X1  g0275(.A1(new_n472), .A2(new_n474), .B1(new_n475), .B2(KEYINPUT6), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n477));
  INV_X1    g0277(.A(G107), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n404), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n307), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n287), .A2(new_n306), .A3(new_n288), .A4(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT83), .B(new_n481), .C1(new_n483), .C2(new_n480), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n479), .A2(new_n285), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n319), .A2(G238), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n346), .B2(new_n319), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n411), .A2(new_n263), .A3(new_n385), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n268), .ZN(new_n495));
  INV_X1    g0295(.A(G45), .ZN(new_n496));
  OAI21_X1  g0296(.A(G250), .B1(new_n496), .B2(G1), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n251), .A2(G45), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n268), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT85), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n257), .B1(new_n492), .B2(new_n493), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n502), .A2(new_n503), .A3(new_n499), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n371), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n500), .ZN(new_n506));
  INV_X1    g0306(.A(G179), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n503), .B1(new_n502), .B2(new_n499), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n307), .A2(new_n353), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G87), .A2(G97), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n478), .B1(new_n260), .B2(new_n207), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n207), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n512), .A2(new_n513), .B1(new_n260), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n411), .A2(new_n207), .A3(new_n263), .A4(new_n385), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n291), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n285), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n353), .B2(new_n483), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n505), .A2(new_n509), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G200), .B1(new_n501), .B2(new_n504), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n506), .A2(G190), .A3(new_n508), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n483), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n467), .A2(G169), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n456), .B(G179), .C1(new_n466), .C2(new_n257), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n488), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n489), .A2(new_n520), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n451), .B1(new_n447), .B2(new_n448), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n455), .A2(G264), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n459), .A2(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n411), .A2(new_n263), .A3(new_n385), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n385), .A2(new_n263), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT90), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n411), .A4(new_n536), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(G257), .A3(G1698), .A4(new_n411), .ZN(new_n542));
  XOR2_X1   g0342(.A(KEYINPUT91), .B(G294), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G33), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n533), .B(new_n535), .C1(new_n545), .C2(new_n268), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G179), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n371), .B2(new_n546), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n478), .A2(KEYINPUT23), .A3(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT23), .B1(new_n478), .B2(G20), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(G20), .B2(new_n493), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n323), .A2(new_n207), .A3(G87), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n552), .A2(new_n523), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(new_n555), .C1(new_n516), .C2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n554), .B1(new_n516), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT24), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n559), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(KEYINPUT88), .A3(KEYINPUT24), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n560), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n285), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n300), .A2(G20), .A3(new_n478), .ZN(new_n569));
  XNOR2_X1  g0369(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n570), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n483), .C2(new_n478), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n548), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n255), .A2(G97), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n577), .B2(new_n462), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n207), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n285), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g0381(.A(new_n581), .B(KEYINPUT20), .Z(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n206), .B2(G33), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n308), .A2(new_n583), .B1(new_n579), .B2(new_n307), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n533), .B1(G270), .B2(new_n455), .ZN(new_n586));
  MUX2_X1   g0386(.A(G257), .B(G264), .S(G1698), .Z(new_n587));
  NAND4_X1  g0387(.A1(new_n411), .A2(new_n263), .A3(new_n385), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n266), .A2(G303), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(KEYINPUT86), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n268), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT86), .B1(new_n588), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n363), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n589), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n268), .A3(new_n590), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(new_n313), .A3(new_n586), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n585), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n371), .B1(new_n582), .B2(new_n584), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(new_n601), .A3(KEYINPUT21), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n585), .A2(new_n598), .A3(G179), .A4(new_n586), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT21), .B1(new_n593), .B2(new_n601), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n535), .B1(new_n545), .B2(new_n268), .ZN(new_n607));
  INV_X1    g0407(.A(new_n533), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n313), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G200), .B2(new_n546), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n568), .A3(new_n574), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n532), .A2(new_n576), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n378), .A2(new_n444), .A3(new_n612), .ZN(G372));
  NOR2_X1   g0413(.A1(new_n378), .A2(new_n444), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n488), .B1(new_n527), .B2(new_n528), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n520), .A2(new_n526), .A3(KEYINPUT26), .A4(new_n615), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT92), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n502), .A2(new_n499), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n525), .B(new_n522), .C1(new_n363), .C2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n509), .B(new_n519), .C1(G169), .C2(new_n618), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n615), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n616), .A2(KEYINPUT92), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n604), .A2(new_n605), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n575), .B2(new_n548), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n619), .A2(new_n620), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n615), .B1(new_n488), .B2(new_n469), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n611), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n620), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n614), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n406), .B(new_n398), .C1(new_n438), .C2(new_n392), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n380), .B1(new_n632), .B2(new_n437), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n427), .B1(new_n633), .B2(new_n429), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n408), .A2(KEYINPUT18), .A3(new_n425), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n315), .A2(new_n359), .B1(new_n283), .B2(new_n310), .ZN(new_n637));
  INV_X1    g0437(.A(new_n423), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n339), .B1(new_n376), .B2(new_n375), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n631), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(new_n300), .ZN(new_n642));
  OR3_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .A3(G20), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT27), .B1(new_n642), .B2(G20), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n585), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n625), .B(new_n606), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n575), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n611), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n576), .ZN(new_n653));
  INV_X1    g0453(.A(new_n576), .ZN(new_n654));
  INV_X1    g0454(.A(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n604), .A2(new_n605), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n647), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n653), .A2(new_n660), .B1(new_n654), .B2(new_n655), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n210), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n663), .A2(KEYINPUT93), .A3(G41), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT93), .B1(new_n663), .B2(G41), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G1), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n511), .A2(new_n478), .A3(new_n579), .ZN(new_n668));
  INV_X1    g0468(.A(new_n216), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n667), .A2(new_n668), .B1(new_n669), .B2(new_n666), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n621), .A2(KEYINPUT26), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n520), .A2(new_n526), .A3(new_n622), .A4(new_n615), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(KEYINPUT29), .B(new_n655), .C1(new_n630), .C2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n620), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n611), .A2(new_n627), .A3(new_n628), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n576), .A2(new_n659), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n617), .A2(new_n623), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n647), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n681), .B2(KEYINPUT29), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n501), .A2(new_n504), .A3(new_n467), .ZN(new_n683));
  OAI211_X1 g0483(.A(G179), .B(new_n586), .C1(new_n591), .C2(new_n592), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n685), .A4(new_n607), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n455), .A2(G257), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n608), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n465), .A2(new_n457), .ZN(new_n689));
  INV_X1    g0489(.A(new_n463), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n688), .B1(new_n691), .B2(new_n268), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n692), .A2(G179), .A3(new_n618), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n607), .A2(new_n608), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n593), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n686), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n508), .A3(new_n506), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n545), .A2(new_n268), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n534), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT30), .B1(new_n700), .B2(new_n685), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n647), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT31), .B(new_n647), .C1(new_n696), .C2(new_n701), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n705), .C1(new_n612), .C2(new_n647), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n682), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n671), .B1(new_n709), .B2(G1), .ZN(G364));
  NOR2_X1   g0510(.A1(new_n299), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n667), .B1(G45), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n650), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n649), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n663), .A2(new_n266), .ZN(new_n717));
  XOR2_X1   g0517(.A(G355), .B(KEYINPUT94), .Z(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n579), .B2(new_n663), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n386), .A2(new_n388), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n210), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n247), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n242), .A2(new_n496), .B1(new_n669), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n213), .B1(G20), .B2(new_n371), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n713), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  NOR4_X1   g0533(.A1(new_n207), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G159), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT97), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n207), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n507), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n266), .B1(new_n745), .B2(G77), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n507), .A2(new_n363), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n742), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n207), .A2(new_n313), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n363), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n746), .B1(new_n291), .B2(new_n748), .C1(new_n523), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n743), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G50), .A2(new_n754), .B1(new_n756), .B2(G58), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n742), .A2(new_n750), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n478), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n207), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n480), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n752), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n741), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(KEYINPUT32), .B2(new_n740), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n737), .B(KEYINPUT98), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(new_n758), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G283), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n266), .B1(new_n755), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n753), .A2(new_n772), .B1(new_n744), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n761), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n771), .B(new_n774), .C1(new_n543), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n748), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  INV_X1    g0578(.A(new_n751), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(G303), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n767), .A2(new_n769), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n765), .A2(KEYINPUT99), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n731), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT99), .B1(new_n765), .B2(new_n781), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n733), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n730), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n649), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n716), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  AOI21_X1  g0590(.A(new_n365), .B1(new_n361), .B2(new_n647), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n359), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n360), .A2(new_n647), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n681), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n655), .B(new_n794), .C1(new_n624), .C2(new_n630), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n707), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n712), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n731), .A2(new_n728), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n712), .B1(G77), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n748), .B1(new_n755), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G303), .B2(new_n754), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n751), .A2(new_n478), .B1(new_n744), .B2(new_n579), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n266), .B1(new_n758), .B2(new_n523), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(new_n762), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n766), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n811), .C1(new_n812), .C2(new_n773), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n720), .B1(new_n394), .B2(new_n761), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n756), .B1(new_n777), .B2(G150), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n754), .A2(G137), .B1(new_n745), .B2(G159), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n751), .A2(new_n202), .B1(new_n758), .B2(new_n291), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT100), .Z(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n813), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n804), .B1(new_n823), .B2(new_n731), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT101), .Z(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n729), .B2(new_n794), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n801), .A2(new_n826), .ZN(G384));
  OAI211_X1 g0627(.A(G116), .B(new_n214), .C1(new_n476), .C2(KEYINPUT35), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(KEYINPUT35), .B2(new_n476), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT36), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n216), .B(G77), .C1(new_n394), .C2(new_n291), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n202), .A2(G68), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n206), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n310), .A2(new_n647), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n311), .A2(new_n315), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n835), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n283), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n283), .A2(KEYINPUT102), .A3(new_n837), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n794), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT30), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n683), .A2(new_n607), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n684), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n686), .A3(new_n695), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT31), .B1(new_n847), .B2(new_n647), .ZN(new_n848));
  INV_X1    g0648(.A(new_n612), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n655), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT105), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n705), .B(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n843), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n400), .A2(new_n289), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n439), .A2(KEYINPUT16), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n380), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n645), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n429), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n408), .A2(new_n420), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n633), .A2(new_n429), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n858), .B1(new_n440), .B2(new_n381), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n860), .A4(new_n854), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n857), .A2(new_n858), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n444), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n869), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n400), .A2(new_n407), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n875), .A2(new_n420), .A3(new_n380), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n425), .B1(new_n875), .B2(new_n380), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT103), .A3(new_n854), .A4(new_n864), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n865), .A2(new_n866), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n879), .A2(new_n880), .B1(KEYINPUT37), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n864), .B1(new_n636), .B2(new_n423), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n853), .A2(new_n885), .A3(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n853), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT81), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n634), .B2(new_n635), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n426), .A2(new_n441), .A3(KEYINPUT81), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n870), .B1(new_n892), .B2(new_n423), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(new_n874), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n869), .B2(new_n872), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT104), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n874), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n873), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n888), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n887), .B1(new_n901), .B2(KEYINPUT40), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n704), .B1(new_n612), .B2(new_n647), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n705), .B(KEYINPUT105), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n614), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n902), .B(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(G330), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n842), .ZN(new_n909));
  INV_X1    g0709(.A(new_n793), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n796), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n898), .A2(new_n899), .A3(new_n873), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n899), .B1(new_n898), .B2(new_n873), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n311), .A2(new_n647), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n873), .A2(new_n884), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n898), .B2(new_n873), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n636), .A2(new_n858), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n675), .B(new_n614), .C1(new_n681), .C2(KEYINPUT29), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n640), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  OAI22_X1  g0725(.A1(new_n908), .A2(new_n925), .B1(new_n206), .B2(new_n711), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n908), .A2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n834), .B1(new_n926), .B2(new_n927), .ZN(G367));
  NAND2_X1  g0728(.A1(new_n711), .A2(G45), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G1), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n628), .B1(new_n488), .B2(new_n655), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n615), .A2(new_n647), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n661), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT44), .B1(new_n661), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n661), .A2(new_n934), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n658), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n650), .A2(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n650), .A2(KEYINPUT109), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n653), .A2(new_n656), .A3(new_n660), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n660), .B1(new_n653), .B2(new_n656), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n945), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(KEYINPUT109), .A3(new_n650), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n709), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n944), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n943), .A2(new_n658), .A3(new_n936), .A4(new_n935), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT110), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n938), .A2(new_n958), .A3(new_n658), .A4(new_n943), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n708), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n666), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n931), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  INV_X1    g0765(.A(new_n934), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n947), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n947), .A2(new_n965), .A3(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT42), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n969), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n967), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n531), .B1(new_n932), .B2(new_n576), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n655), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n525), .A2(new_n655), .ZN(new_n977));
  MUX2_X1   g0777(.A(new_n627), .B(new_n676), .S(new_n977), .Z(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT43), .Z(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(KEYINPUT108), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT108), .B1(new_n976), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n970), .A2(new_n973), .A3(new_n975), .A4(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT107), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n983), .A2(new_n987), .B1(new_n658), .B2(new_n966), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n985), .B(KEYINPUT107), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n658), .A2(new_n966), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n982), .C2(new_n981), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n964), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n732), .B1(new_n210), .B2(new_n353), .C1(new_n724), .C2(new_n238), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(new_n712), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G143), .A2(new_n754), .B1(new_n756), .B2(G150), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n291), .B2(new_n761), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT112), .Z(new_n997));
  OAI22_X1  g0797(.A1(new_n748), .A2(new_n738), .B1(new_n758), .B2(new_n293), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G50), .B2(new_n745), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n266), .B1(new_n779), .B2(G58), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT113), .B(G137), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1000), .C1(new_n737), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n737), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(G317), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n543), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1005), .A2(new_n748), .B1(new_n773), .B2(new_n753), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G283), .B2(new_n745), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n758), .A2(new_n480), .ZN(new_n1008));
  INV_X1    g0808(.A(G303), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n755), .A2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G107), .C2(new_n775), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT46), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n751), .B2(new_n579), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1004), .A2(new_n1007), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n779), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n721), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n997), .A2(new_n1002), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT114), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n731), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n994), .B1(new_n787), .B2(new_n978), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n992), .A2(new_n1024), .ZN(G387));
  AOI21_X1  g0825(.A(new_n931), .B1(new_n950), .B2(new_n952), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT115), .Z(new_n1027));
  OAI22_X1  g0827(.A1(new_n748), .A2(new_n331), .B1(new_n744), .B2(new_n291), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT116), .Z(new_n1029));
  NAND2_X1  g0829(.A1(new_n1003), .A2(G150), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n753), .A2(new_n738), .B1(new_n755), .B2(new_n202), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n761), .A2(new_n353), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n751), .A2(new_n293), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1008), .A4(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n720), .A3(new_n1030), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n744), .A2(new_n1009), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n773), .A2(new_n748), .B1(new_n755), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1036), .B(new_n1038), .C1(G322), .C2(new_n754), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT48), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(KEYINPUT48), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n775), .A2(G283), .B1(new_n779), .B2(new_n543), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT49), .Z(new_n1044));
  OAI221_X1 g0844(.A(new_n721), .B1(new_n579), .B2(new_n758), .C1(new_n737), .C2(new_n772), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1035), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT117), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(KEYINPUT117), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n731), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n657), .A2(new_n730), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n724), .B1(new_n234), .B2(new_n725), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n668), .B2(new_n717), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n351), .B2(new_n202), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n331), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n496), .B1(new_n291), .B2(new_n293), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n668), .A4(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1052), .A2(new_n1057), .B1(G107), .B2(new_n210), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n713), .B1(new_n1058), .B2(new_n732), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1049), .A2(new_n1050), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n709), .A2(new_n953), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT118), .B2(new_n954), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n666), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1027), .B(new_n1060), .C1(new_n1062), .C2(new_n1065), .ZN(G393));
  OAI221_X1 g0866(.A(new_n732), .B1(new_n480), .B2(new_n210), .C1(new_n724), .C2(new_n245), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(new_n712), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n777), .B1(new_n779), .B2(G68), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G87), .A2(new_n768), .B1(new_n745), .B2(new_n351), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n775), .A2(G77), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(G150), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n753), .A2(new_n1073), .B1(new_n755), .B2(new_n738), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1003), .A2(G143), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1075), .A3(new_n1076), .A4(new_n720), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n748), .A2(new_n1009), .B1(new_n744), .B2(new_n806), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n266), .B1(new_n758), .B2(new_n478), .C1(new_n761), .C2(new_n579), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G283), .C2(new_n779), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n753), .A2(new_n1037), .B1(new_n755), .B2(new_n773), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT121), .Z(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT120), .B(KEYINPUT52), .Z(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1080), .B1(new_n770), .B2(new_n737), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1082), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1077), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT122), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n731), .B1(new_n1088), .B2(KEYINPUT122), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1068), .B1(new_n1089), .B2(new_n1090), .C1(new_n934), .C2(new_n787), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT119), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n937), .B1(new_n942), .B2(new_n941), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n658), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n944), .A2(KEYINPUT119), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n960), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1096), .B2(new_n931), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n954), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n666), .B1(new_n955), .B2(new_n960), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  AOI21_X1  g0901(.A(new_n915), .B1(new_n873), .B2(new_n884), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n674), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n647), .B1(new_n679), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n792), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n793), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1102), .B1(new_n1106), .B2(new_n909), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n706), .A2(G330), .A3(new_n794), .A4(new_n842), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT39), .B1(new_n895), .B2(new_n896), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(KEYINPUT39), .B2(new_n885), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n796), .A2(new_n910), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n915), .B1(new_n1111), .B2(new_n842), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1107), .B(new_n1108), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n793), .B1(new_n681), .B2(new_n794), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1114), .A2(new_n909), .B1(new_n311), .B2(new_n647), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n917), .A2(new_n918), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n655), .B(new_n1105), .C1(new_n630), .C2(new_n674), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n842), .B1(new_n1118), .B2(new_n793), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1115), .A2(new_n1116), .B1(new_n1119), .B2(new_n1102), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n794), .A2(G330), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n842), .C1(new_n904), .C2(new_n903), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1113), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1116), .A2(new_n728), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n712), .B1(new_n351), .B2(new_n803), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n812), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n779), .A2(G150), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n755), .A2(new_n814), .B1(new_n758), .B2(new_n202), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n753), .A2(new_n1133), .B1(new_n748), .B2(new_n1001), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n323), .B1(new_n744), .B2(new_n1135), .C1(new_n761), .C2(new_n738), .ZN(new_n1136));
  OR4_X1    g0936(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n812), .A2(new_n806), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n753), .A2(new_n805), .B1(new_n748), .B2(new_n478), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G97), .B2(new_n745), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n323), .B1(new_n779), .B2(G87), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G116), .A2(new_n756), .B1(new_n768), .B2(G68), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n1071), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1129), .A2(new_n1137), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1127), .B1(new_n1144), .B2(new_n731), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1125), .A2(new_n930), .B1(new_n1126), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n614), .B(G330), .C1(new_n904), .C2(new_n903), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n923), .A2(new_n1147), .A3(new_n640), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n706), .A2(G330), .A3(new_n794), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n909), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1123), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1111), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1121), .B1(new_n850), .B2(new_n852), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1106), .B(new_n1108), .C1(new_n842), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n1113), .C1(new_n1120), .C2(new_n1123), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(KEYINPUT123), .A3(new_n1064), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1124), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT123), .B1(new_n1156), .B2(new_n1064), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1146), .B1(new_n1160), .B2(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n339), .A2(new_n373), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(new_n336), .A3(new_n858), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n336), .A2(new_n858), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n339), .A2(new_n373), .A3(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1164), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n922), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n887), .B(G330), .C1(new_n901), .C2(KEYINPUT40), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n914), .A2(new_n919), .A3(new_n1171), .A4(new_n921), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n930), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n758), .A2(new_n394), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n720), .A2(G41), .A3(new_n1033), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n812), .B2(new_n805), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT124), .Z(new_n1182));
  OAI22_X1  g0982(.A1(new_n748), .A2(new_n480), .B1(new_n744), .B2(new_n353), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n753), .A2(new_n579), .B1(new_n755), .B2(new_n478), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G68), .C2(new_n775), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n255), .B(new_n248), .C1(new_n758), .C2(new_n738), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1003), .A2(G124), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n753), .A2(new_n1128), .B1(new_n748), .B2(new_n814), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G150), .B2(new_n775), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n745), .A2(G137), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1135), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1194), .A2(new_n779), .B1(new_n756), .B2(G128), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1189), .B(new_n1190), .C1(KEYINPUT59), .C2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n248), .B1(new_n721), .B2(new_n255), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1197), .A2(new_n1198), .B1(new_n202), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1187), .B2(KEYINPUT58), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n731), .B1(new_n1188), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n713), .B1(new_n202), .B2(new_n802), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n1172), .C2(new_n729), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1178), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1148), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1156), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n853), .B1(new_n912), .B2(new_n913), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT40), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n907), .B(new_n886), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n897), .A2(new_n900), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n920), .B1(new_n1213), .B2(new_n911), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1171), .B1(new_n1214), .B2(new_n919), .ZN(new_n1215));
  AND4_X1   g1015(.A1(new_n919), .A2(new_n914), .A3(new_n921), .A4(new_n1171), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1212), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT57), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1207), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1209), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1205), .B1(new_n1222), .B2(new_n1064), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1153), .A2(new_n842), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1114), .B1(new_n1123), .B2(new_n1150), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n930), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(KEYINPUT125), .A3(new_n930), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n909), .A2(new_n728), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n712), .B1(G68), .B2(new_n803), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n812), .A2(new_n1009), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n755), .A2(new_n805), .B1(new_n744), .B2(new_n478), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G294), .B2(new_n754), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1032), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n323), .B1(new_n768), .B2(G77), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G97), .A2(new_n779), .B1(new_n777), .B2(G116), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n812), .A2(new_n1133), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n753), .A2(new_n814), .B1(new_n755), .B2(new_n1001), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n748), .A2(new_n1135), .B1(new_n744), .B2(new_n1073), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n775), .A2(G50), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1179), .B1(G159), .B2(new_n779), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n720), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1236), .A2(new_n1242), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1235), .B1(new_n1250), .B2(new_n731), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1231), .A2(new_n1233), .B1(new_n1234), .B2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1148), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n962), .A3(new_n1158), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(G381));
  NOR2_X1   g1056(.A1(G375), .A2(G378), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1100), .A2(new_n992), .A3(new_n1024), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(G407));
  INV_X1    g1061(.A(G213), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G343), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  XNOR2_X1  g1065(.A(G393), .B(new_n789), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1100), .B1(new_n992), .B2(new_n1024), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1259), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(G390), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1266), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1258), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1155), .A2(new_n666), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1253), .B2(new_n1148), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1232), .A2(KEYINPUT60), .A3(new_n1206), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1252), .A3(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1252), .A3(new_n1280), .A4(G384), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1252), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1279), .A2(new_n1281), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1263), .ZN(new_n1286));
  INV_X1    g1086(.A(G2897), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1279), .A2(new_n1281), .A3(new_n1284), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1287), .B2(new_n1286), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1178), .A2(new_n1204), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1219), .A2(new_n962), .A3(new_n1207), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1223), .B2(G378), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(new_n1263), .ZN(new_n1297));
  AOI221_X4 g1097(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1206), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1220), .B1(new_n1219), .B2(new_n1207), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1064), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G378), .A3(new_n1293), .ZN(new_n1301));
  INV_X1    g1101(.A(G378), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(new_n1178), .A3(new_n1204), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1286), .A4(new_n1285), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1297), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1263), .B(new_n1290), .C1(new_n1301), .C2(new_n1304), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(new_n1306), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1272), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1305), .A2(new_n1286), .A3(new_n1285), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1305), .A2(new_n1286), .B1(new_n1291), .B2(new_n1289), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1268), .A2(new_n1271), .A3(new_n1308), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(KEYINPUT63), .B2(new_n1310), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1312), .A2(new_n1319), .A3(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(G405));
  XNOR2_X1  g1124(.A(new_n1223), .B(G378), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1272), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1285), .ZN(G402));
endmodule


