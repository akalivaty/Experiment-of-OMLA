//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n208), .B(new_n214), .C1(G58), .C2(G232), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n207), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT86), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  OAI211_X1 g0045(.A(G1), .B(G13), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT64), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n244), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT84), .B(G303), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n213), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(G264), .C2(new_n258), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n246), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT5), .A2(G41), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT5), .A2(G41), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n263), .B(G274), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n265), .B2(new_n264), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n268), .A2(G270), .A3(new_n246), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n261), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G200), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT65), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(new_n220), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n273), .B2(new_n220), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G116), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n206), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G283), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(new_n219), .C1(G33), .C2(new_n212), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n273), .A2(new_n220), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n206), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT20), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(new_n284), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n243), .B1(new_n272), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n270), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(new_n294), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(KEYINPUT86), .C1(new_n270), .C2(new_n271), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n269), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n256), .A2(new_n260), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n266), .B(new_n300), .C1(new_n301), .C2(new_n246), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT21), .A3(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n270), .A2(G179), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n294), .A3(G169), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT21), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT85), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(KEYINPUT85), .A3(new_n308), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n299), .A2(new_n306), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT19), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n219), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G97), .A2(G107), .ZN(new_n317));
  INV_X1    g0117(.A(G87), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n219), .B(G68), .C1(new_n247), .C2(new_n248), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n315), .B1(new_n314), .B2(G20), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n287), .A2(KEYINPUT65), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n275), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n279), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT82), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n324), .A2(new_n278), .A3(new_n275), .A4(new_n282), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n281), .A2(KEYINPUT82), .A3(G87), .A4(new_n282), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(G244), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT81), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n257), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n257), .A2(G238), .A3(new_n258), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G116), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n246), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n263), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G250), .B1(G274), .B2(new_n263), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT70), .B(G200), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT83), .B(new_n335), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT83), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n334), .A2(new_n333), .ZN(new_n352));
  INV_X1    g0152(.A(new_n330), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n344), .B2(new_n346), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(G190), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n350), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n344), .A2(new_n346), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n281), .A2(new_n327), .A3(new_n282), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT68), .B(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n347), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n313), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G20), .A2(G33), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT6), .ZN(new_n373));
  INV_X1    g0173(.A(G107), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n212), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n375), .B2(new_n317), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(KEYINPUT6), .A3(G97), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n219), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n249), .A2(new_n254), .A3(new_n219), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n247), .A2(new_n248), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n372), .B(new_n380), .C1(new_n389), .C2(new_n374), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n325), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n249), .A2(new_n254), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G250), .A3(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT4), .ZN(new_n394));
  INV_X1    g0194(.A(G244), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT64), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n258), .B(new_n396), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n257), .A2(G244), .A3(new_n258), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n394), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n393), .A2(new_n399), .A3(new_n401), .A4(new_n285), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n343), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n268), .A2(G257), .A3(new_n246), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT78), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n404), .A2(new_n405), .A3(new_n266), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n404), .B2(new_n266), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n266), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n402), .B2(new_n343), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n409), .A2(G200), .B1(new_n411), .B2(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n332), .A2(G97), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G97), .B2(new_n279), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND4_X1   g0217(.A1(KEYINPUT79), .A2(new_n391), .A3(new_n412), .A4(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n390), .A2(new_n325), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT79), .B1(new_n419), .B2(new_n412), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n381), .A2(new_n383), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n387), .A3(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n371), .B(new_n379), .C1(new_n425), .C2(G107), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n276), .A2(new_n280), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n417), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n411), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n360), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n403), .A2(new_n363), .A3(new_n408), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n403), .A2(KEYINPUT80), .A3(new_n363), .A4(new_n408), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n428), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT23), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n219), .B2(G107), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n374), .A2(KEYINPUT23), .A3(G20), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n244), .A2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(new_n439), .B1(new_n440), .B2(G116), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT22), .A2(G20), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n392), .A2(G87), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n257), .A2(new_n219), .A3(G87), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT22), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n443), .A2(KEYINPUT87), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT87), .B1(new_n443), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT24), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(KEYINPUT24), .B(new_n441), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n325), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT25), .B1(new_n278), .B2(G107), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n278), .A2(KEYINPUT25), .A3(G107), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n332), .C2(new_n374), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT88), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT89), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G294), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n257), .A2(G250), .A3(new_n258), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT89), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n257), .A2(new_n461), .A3(G257), .A4(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n343), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n268), .A2(new_n246), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT90), .A3(G264), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n268), .A2(G264), .A3(new_n246), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT90), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n464), .A2(new_n266), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n271), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n463), .A2(new_n343), .B1(new_n466), .B2(new_n469), .ZN(new_n473));
  INV_X1    g0273(.A(G190), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n266), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n452), .A2(new_n456), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n360), .ZN(new_n478));
  INV_X1    g0278(.A(G179), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n473), .A2(new_n479), .A3(new_n266), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n452), .B2(new_n456), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n367), .A2(new_n421), .A3(new_n436), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT13), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n392), .A2(G232), .A3(G1698), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT72), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n487), .A2(new_n392), .A3(G226), .A4(new_n258), .ZN(new_n488));
  AOI21_X1  g0288(.A(G1698), .B1(new_n249), .B2(new_n254), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(G226), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n314), .B(new_n486), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n343), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n246), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n211), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G274), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n485), .A2(new_n492), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n491), .B2(new_n343), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n485), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT14), .ZN(new_n504));
  INV_X1    g0304(.A(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(G179), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT14), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(G169), .C1(new_n500), .C2(new_n502), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n277), .A2(G20), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n427), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT12), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n279), .A2(new_n210), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n513), .A2(G68), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n440), .A2(G77), .B1(new_n368), .B2(G50), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n219), .B2(G68), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n325), .ZN(new_n520));
  XOR2_X1   g0320(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT11), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n520), .B(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n510), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT8), .B(G58), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n368), .B1(new_n327), .B2(new_n440), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n219), .B2(new_n370), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n325), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n513), .A2(G77), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n279), .A2(new_n370), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n392), .A2(G238), .A3(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n374), .B2(new_n392), .ZN(new_n536));
  INV_X1    g0336(.A(new_n392), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n537), .A2(new_n228), .A3(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n343), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n499), .B1(new_n494), .B2(new_n395), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT69), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n534), .B1(new_n543), .B2(new_n363), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n360), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n257), .B1(G223), .B2(G1698), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n258), .A2(G226), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n548), .A2(new_n549), .B1(new_n244), .B2(new_n318), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n498), .B1(new_n550), .B2(new_n343), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n494), .A2(new_n228), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n363), .A3(new_n553), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n498), .B(new_n552), .C1(new_n550), .C2(new_n343), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G159), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n369), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g0359(.A(KEYINPUT66), .B(G58), .Z(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G68), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n202), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(G20), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n383), .B1(new_n257), .B2(G20), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n210), .B1(new_n564), .B2(new_n387), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT16), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n325), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n563), .B1(new_n389), .B2(new_n210), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n568), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT8), .ZN(new_n572));
  OR2_X1    g0372(.A1(KEYINPUT66), .A2(G58), .ZN(new_n573));
  NAND2_X1  g0373(.A1(KEYINPUT66), .A2(G58), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n572), .A2(G58), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n279), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n512), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n557), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT18), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n201), .B1(new_n560), .B2(G68), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n583), .A2(new_n219), .B1(new_n558), .B2(new_n369), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n565), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n427), .B1(new_n585), .B2(KEYINPUT16), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n425), .B2(G68), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT16), .ZN(new_n588));
  INV_X1    g0388(.A(new_n579), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n556), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n555), .A2(new_n474), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n555), .B2(G200), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT17), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT17), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n588), .A2(new_n593), .A3(new_n596), .A4(new_n589), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n582), .A2(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n542), .A2(new_n348), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(new_n534), .C1(new_n474), .C2(new_n542), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n392), .A2(G223), .A3(G1698), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n392), .A2(G222), .A3(new_n258), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n249), .A2(new_n254), .A3(G77), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n343), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n246), .A2(G226), .A3(new_n493), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n499), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n360), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n278), .A2(G50), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n440), .B1(new_n575), .B2(new_n576), .ZN(new_n610));
  INV_X1    g0410(.A(G50), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n219), .B1(new_n201), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT67), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n368), .A2(G150), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(KEYINPUT67), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n610), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n609), .B1(new_n616), .B2(new_n325), .ZN(new_n617));
  AND4_X1   g0417(.A1(G50), .A2(new_n324), .A3(new_n511), .A4(new_n275), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g0420(.A(KEYINPUT68), .B(G179), .Z(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n607), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT71), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT9), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n624), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n609), .B(new_n618), .C1(new_n616), .C2(new_n325), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(KEYINPUT9), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n607), .A2(new_n348), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n605), .A2(G190), .A3(new_n499), .A4(new_n606), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT71), .B1(new_n627), .B2(KEYINPUT9), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n620), .A2(new_n625), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n631), .A3(new_n635), .A4(new_n632), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT10), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n623), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n505), .A2(G190), .A3(new_n506), .ZN(new_n639));
  OAI21_X1  g0439(.A(G200), .B1(new_n500), .B2(new_n502), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(new_n524), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n598), .A2(new_n600), .A3(new_n638), .A4(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT76), .B1(new_n547), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n598), .A2(new_n638), .A3(new_n641), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n510), .A2(new_n525), .B1(new_n545), .B2(new_n544), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT76), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .A4(new_n600), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n484), .B1(new_n643), .B2(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n595), .A2(new_n597), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n547), .A2(new_n649), .A3(new_n641), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n588), .A2(new_n589), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT18), .B1(new_n652), .B2(new_n557), .ZN(new_n653));
  AOI211_X1 g0453(.A(new_n581), .B(new_n556), .C1(new_n588), .C2(new_n589), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n582), .A2(KEYINPUT91), .A3(new_n591), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n637), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n623), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n643), .A2(new_n647), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n436), .B2(new_n366), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n391), .A2(new_n417), .B1(new_n433), .B2(new_n434), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n354), .A2(new_n355), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n357), .A2(new_n668), .B1(new_n362), .B2(new_n364), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n430), .A4(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n665), .A2(new_n365), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n452), .A2(new_n456), .ZN(new_n673));
  INV_X1    g0473(.A(new_n481), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n312), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT85), .B1(new_n307), .B2(new_n308), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n676), .A2(new_n305), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n452), .A2(new_n456), .A3(new_n476), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n421), .A3(new_n436), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n663), .B1(new_n664), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT92), .ZN(G369));
  NAND3_X1  g0484(.A1(new_n306), .A2(new_n311), .A3(new_n312), .ZN(new_n685));
  INV_X1    g0485(.A(G13), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G20), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n277), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n297), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n313), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT93), .B(G330), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n673), .A2(new_n693), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n483), .A2(new_n700), .B1(new_n482), .B2(new_n693), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AND4_X1   g0503(.A1(new_n483), .A2(new_n685), .A3(new_n694), .A4(new_n700), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n675), .A2(new_n693), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n223), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n319), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n710), .A2(new_n218), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(KEYINPUT94), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(KEYINPUT94), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n411), .A2(new_n473), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n304), .A3(new_n359), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n270), .A2(new_n621), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n409), .A3(new_n471), .A4(new_n359), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n693), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT31), .B(new_n724), .C1(new_n484), .C2(new_n693), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n698), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n428), .A2(new_n430), .A3(new_n435), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n358), .A2(new_n365), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n667), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n436), .B2(new_n672), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n365), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n391), .A2(new_n412), .A3(new_n417), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT79), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n419), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(new_n436), .A3(new_n737), .A4(new_n680), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n669), .B1(new_n685), .B2(new_n482), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n694), .C1(new_n733), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n693), .B1(new_n671), .B2(new_n681), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n742), .B2(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n716), .B1(new_n745), .B2(G1), .ZN(G364));
  NAND2_X1  g0546(.A1(new_n687), .A2(G45), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n710), .A2(G1), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n697), .B2(new_n698), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n698), .B2(new_n697), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n220), .B1(G20), .B2(new_n360), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n218), .A2(G45), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n238), .B2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n708), .A2(new_n257), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n759), .A2(new_n760), .B1(new_n206), .B2(new_n708), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n392), .A2(G355), .A3(new_n223), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n474), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n219), .B1(new_n764), .B2(new_n479), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G97), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n219), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n348), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n474), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G87), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  AND4_X1   g0574(.A1(new_n392), .A2(new_n768), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n621), .A2(KEYINPUT95), .A3(G20), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT95), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n363), .B2(new_n219), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n474), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(G190), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G50), .A2(new_n781), .B1(new_n782), .B2(G68), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n764), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n560), .A2(new_n785), .B1(new_n787), .B2(G77), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n769), .A2(new_n786), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n558), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n775), .A2(new_n783), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n789), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G329), .ZN(new_n794));
  INV_X1    g0594(.A(new_n773), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n771), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n537), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n797), .B(new_n801), .C1(G326), .C2(new_n781), .ZN(new_n802));
  INV_X1    g0602(.A(new_n782), .ZN(new_n803));
  INV_X1    g0603(.A(G317), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(KEYINPUT33), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(KEYINPUT33), .B2(new_n804), .ZN(new_n806));
  INV_X1    g0606(.A(new_n787), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n807), .A2(new_n808), .B1(KEYINPUT97), .B2(new_n800), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G322), .B2(new_n785), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n802), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n765), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n792), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n763), .B1(new_n814), .B2(new_n755), .ZN(new_n815));
  INV_X1    g0615(.A(new_n754), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n749), .C1(new_n697), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n751), .A2(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n546), .A2(new_n693), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n600), .B1(new_n534), .B2(new_n694), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n546), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n742), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n748), .B1(new_n728), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n728), .A2(new_n822), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(KEYINPUT102), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n825), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n781), .A2(G137), .B1(G159), .B2(new_n787), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n784), .C1(new_n833), .C2(new_n803), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT34), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n795), .A2(new_n210), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n257), .B1(new_n789), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n771), .A2(G50), .B1(new_n838), .B2(KEYINPUT99), .ZN(new_n839));
  INV_X1    g0639(.A(new_n560), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(KEYINPUT99), .B2(new_n838), .C1(new_n840), .C2(new_n765), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n785), .A2(G294), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n537), .B1(new_n808), .B2(new_n789), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G87), .B2(new_n773), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n771), .A2(G107), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n768), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n781), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT98), .B(G283), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n799), .A2(new_n848), .B1(new_n803), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n847), .B(new_n851), .C1(G116), .C2(new_n787), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n755), .B1(new_n842), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n755), .A2(new_n752), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n370), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n749), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT100), .Z(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n753), .B2(new_n821), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n830), .A2(new_n858), .ZN(G384));
  INV_X1    g0659(.A(new_n691), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n658), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n585), .A2(KEYINPUT16), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n589), .B1(new_n569), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n557), .B2(new_n860), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n865), .B2(new_n594), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n652), .A2(new_n860), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n867), .A2(new_n580), .A3(new_n594), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n866), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n864), .A2(new_n860), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n598), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n594), .A2(KEYINPUT17), .ZN(new_n874));
  INV_X1    g0674(.A(new_n597), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n874), .A2(new_n875), .B1(new_n653), .B2(new_n654), .ZN(new_n876));
  INV_X1    g0676(.A(new_n872), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT104), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n870), .B(KEYINPUT38), .C1(new_n873), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n867), .A2(new_n580), .A3(new_n594), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n862), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n691), .B1(new_n588), .B2(new_n589), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n655), .A2(new_n656), .A3(new_n649), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n879), .B(new_n880), .C1(new_n885), .C2(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT105), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n871), .B1(new_n598), .B2(new_n872), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n876), .A2(KEYINPUT104), .A3(new_n877), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n890), .B2(new_n870), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n892), .B(new_n869), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT39), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n884), .A2(new_n883), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n880), .A4(new_n879), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n887), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n510), .A2(new_n525), .A3(new_n694), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n861), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n891), .A2(new_n893), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n665), .A2(new_n365), .A3(new_n670), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n821), .B(new_n694), .C1(new_n740), .C2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n546), .B2(new_n693), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n525), .A2(new_n693), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n526), .A2(new_n641), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n641), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n525), .B(new_n693), .C1(new_n909), .C2(new_n510), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT107), .Z(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n911), .A2(new_n725), .A3(new_n726), .A4(new_n821), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n903), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n908), .A2(new_n910), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n725), .A2(new_n726), .A3(new_n821), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n896), .A2(new_n879), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n664), .A2(new_n727), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n924), .B(new_n925), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n698), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n915), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n743), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n664), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n664), .A3(KEYINPUT106), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n663), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n928), .B(new_n934), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n277), .B2(new_n687), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT35), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n219), .B(new_n220), .C1(new_n378), .C2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(G116), .C1(new_n937), .C2(new_n378), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT103), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n561), .A2(G50), .A3(G77), .A4(new_n202), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(G50), .B2(new_n210), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n686), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(new_n941), .A3(new_n944), .ZN(G367));
  AOI21_X1  g0745(.A(KEYINPUT46), .B1(new_n771), .B2(G116), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n257), .B(new_n946), .C1(G317), .C2(new_n793), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n773), .A2(G97), .ZN(new_n949));
  INV_X1    g0749(.A(new_n765), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(G107), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n787), .B2(new_n849), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n785), .A2(new_n255), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT113), .B(G311), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G294), .A2(new_n782), .B1(new_n781), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n803), .A2(new_n558), .B1(new_n807), .B2(new_n611), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n766), .A2(new_n210), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G150), .B2(new_n785), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n795), .A2(new_n370), .ZN(new_n963));
  INV_X1    g0763(.A(G137), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n392), .B1(new_n964), .B2(new_n789), .C1(new_n798), .C2(new_n840), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(new_n781), .C2(G143), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n960), .A3(new_n962), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n957), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT115), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n755), .ZN(new_n971));
  INV_X1    g0771(.A(new_n760), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n756), .B1(new_n223), .B2(new_n328), .C1(new_n234), .C2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n335), .A2(new_n694), .ZN(new_n974));
  MUX2_X1   g0774(.A(new_n672), .B(new_n365), .S(new_n974), .Z(new_n975));
  AOI21_X1  g0775(.A(new_n748), .B1(new_n975), .B2(new_n754), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n975), .B(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n428), .A2(new_n693), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n736), .A2(new_n436), .A3(new_n737), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n729), .A2(new_n693), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT108), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT108), .B1(new_n981), .B2(new_n982), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n436), .B1(new_n987), .B2(new_n675), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n983), .B(new_n984), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n704), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n988), .A2(new_n694), .B1(new_n990), .B2(KEYINPUT42), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT42), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n704), .C1(new_n985), .C2(new_n986), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT109), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n996), .B1(new_n991), .B2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n979), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n991), .A2(new_n995), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT110), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n975), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1004), .A3(new_n997), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n987), .A2(new_n703), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n978), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1000), .A2(new_n1005), .A3(KEYINPUT111), .A4(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n747), .A2(G1), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n706), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT112), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT44), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1016), .A2(new_n987), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n989), .C2(new_n706), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n989), .A2(KEYINPUT45), .A3(new_n706), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT45), .B1(new_n989), .B2(new_n706), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1019), .B(new_n1022), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n702), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n685), .A2(new_n694), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n704), .B1(new_n701), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(new_n699), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n744), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1016), .B2(new_n987), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n1023), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1034), .A2(new_n703), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1027), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1015), .B1(new_n1036), .B2(new_n745), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1012), .B1(new_n1013), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n977), .B1(new_n1011), .B2(new_n1038), .ZN(G387));
  OAI21_X1  g0839(.A(new_n386), .B1(new_n795), .B2(new_n206), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n781), .A2(G322), .B1(new_n255), .B2(new_n787), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n782), .A2(new_n955), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n804), .C2(new_n784), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT48), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n812), .B2(new_n798), .C1(new_n765), .C2(new_n850), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT49), .Z(new_n1046));
  AOI211_X1 g0846(.A(new_n1040), .B(new_n1046), .C1(G326), .C2(new_n793), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n803), .A2(new_n577), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G50), .A2(new_n785), .B1(new_n787), .B2(G68), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n767), .A2(new_n327), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n257), .B1(new_n789), .B2(new_n833), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n771), .B2(G77), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n949), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1048), .B(new_n1053), .C1(G159), .C2(new_n781), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n755), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n701), .A2(new_n754), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n527), .A2(G50), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT50), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n711), .B1(new_n210), .B2(new_n370), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(G45), .B(new_n1059), .C1(new_n1058), .C2(new_n1057), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n760), .B1(new_n231), .B2(new_n262), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n392), .B(new_n223), .C1(G116), .C2(new_n319), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n223), .A2(G107), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n756), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1055), .A2(new_n749), .A3(new_n1056), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1031), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n710), .B1(new_n744), .B2(new_n1030), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1013), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1066), .B(new_n1069), .C1(new_n1070), .C2(new_n1030), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1067), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n709), .A3(new_n1036), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1027), .A2(new_n1035), .A3(new_n1013), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n223), .A2(new_n212), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n757), .B(new_n1076), .C1(new_n241), .C2(new_n760), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n774), .B1(new_n798), .B2(new_n850), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n392), .B(new_n1078), .C1(G116), .C2(new_n950), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n812), .B2(new_n807), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n255), .B2(new_n782), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n793), .A2(G322), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n781), .A2(G317), .B1(new_n785), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1081), .A2(new_n1082), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n781), .A2(G150), .B1(new_n785), .B2(G159), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT51), .Z(new_n1089));
  NOR2_X1   g0889(.A1(new_n766), .A2(new_n370), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n257), .B1(new_n832), .B2(new_n789), .C1(new_n798), .C2(new_n210), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n782), .C2(G50), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n787), .A2(new_n528), .B1(G87), .B2(new_n773), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n748), .B(new_n1077), .C1(new_n1095), .C2(new_n755), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT117), .Z(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n816), .B2(new_n989), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1074), .A2(new_n1075), .A3(new_n1098), .ZN(G390));
  NAND4_X1  g0899(.A1(new_n725), .A2(G330), .A3(new_n726), .A4(new_n821), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n919), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n725), .A2(new_n698), .A3(new_n726), .A4(new_n821), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n919), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n820), .A2(new_n546), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n694), .B(new_n1105), .C1(new_n733), .C2(new_n740), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n819), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1102), .A2(new_n919), .ZN(new_n1109));
  INV_X1    g0909(.A(G330), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n917), .B2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1104), .A2(new_n1108), .B1(new_n1111), .B2(new_n906), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n623), .B1(new_n659), .B2(new_n660), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n664), .A2(G330), .A3(new_n727), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n664), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT106), .B1(new_n929), .B2(new_n664), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1113), .B(new_n1114), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT118), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1111), .A2(new_n906), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1100), .A2(new_n919), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n1108), .C1(new_n919), .C2(new_n1102), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n934), .A3(new_n1123), .A4(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n912), .A2(new_n900), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n887), .A2(new_n1126), .A3(new_n894), .A4(new_n898), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n922), .B(new_n900), .C1(new_n919), .C2(new_n1108), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1103), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n917), .A2(new_n1110), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n709), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n537), .B1(new_n812), .B2(new_n789), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1090), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n772), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n807), .A2(new_n212), .B1(new_n206), .B2(new_n784), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n836), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n374), .B2(new_n803), .C1(new_n796), .C2(new_n848), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n789), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n392), .B1(new_n795), .B2(new_n611), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n798), .A2(new_n833), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT53), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n558), .B2(new_n766), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1144), .B(new_n1147), .C1(new_n1146), .C2(new_n1145), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G128), .A2(new_n781), .B1(new_n782), .B2(G137), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT54), .B(G143), .Z(new_n1150));
  AOI22_X1  g0950(.A1(G132), .A2(new_n785), .B1(new_n787), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(new_n755), .B1(new_n577), .B2(new_n854), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n749), .B(new_n1154), .C1(new_n899), .C2(new_n753), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1132), .B2(new_n1013), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1135), .A2(new_n1157), .A3(new_n1159), .ZN(G378));
  AOI22_X1  g0960(.A1(new_n785), .A2(G128), .B1(new_n767), .B2(G150), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n964), .B2(new_n807), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1142), .A2(new_n848), .B1(new_n803), .B2(new_n837), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n771), .C2(new_n1150), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT59), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n773), .B2(G159), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT120), .B(G124), .Z(new_n1167));
  AOI21_X1  g0967(.A(G33), .B1(new_n793), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n212), .A2(new_n803), .B1(new_n848), .B2(new_n206), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n386), .B1(new_n796), .B2(new_n789), .C1(new_n795), .C2(new_n840), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n245), .B1(new_n798), .B2(new_n370), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1171), .A2(new_n961), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n328), .B2(new_n807), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1170), .B(new_n1174), .C1(G107), .C2(new_n785), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT58), .Z(new_n1176));
  OAI21_X1  g0976(.A(new_n611), .B1(new_n247), .B2(G41), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n748), .B1(new_n1178), .B2(new_n755), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n627), .A2(new_n691), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n638), .B(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT55), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT56), .ZN(new_n1185));
  OR3_X1    g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1179), .B1(new_n1188), .B2(new_n753), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n611), .B2(new_n854), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n918), .A2(G330), .A3(new_n923), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n918), .A2(new_n1188), .A3(G330), .A4(new_n923), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(new_n914), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n1196), .B2(new_n1013), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1117), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1134), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1196), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n913), .A2(new_n1193), .A3(new_n902), .A4(new_n1194), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1194), .A2(new_n1193), .B1(new_n902), .B2(new_n913), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1117), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n709), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1197), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1197), .C1(new_n1200), .C2(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n919), .A2(new_n752), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n766), .A2(new_n611), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n386), .B(new_n1212), .C1(G128), .C2(new_n793), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G159), .A2(new_n771), .B1(new_n773), .B2(new_n560), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n833), .C2(new_n807), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n782), .B2(new_n1150), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n781), .A2(G132), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT123), .Z(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n964), .C2(new_n784), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1050), .B1(new_n784), .B2(new_n796), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  OAI221_X1 g1021(.A(new_n537), .B1(new_n799), .B2(new_n789), .C1(new_n807), .C2(new_n374), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G294), .B2(new_n781), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n798), .A2(new_n212), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n963), .B(new_n1224), .C1(new_n782), .C2(G116), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1227), .A2(new_n755), .B1(new_n210), .B2(new_n854), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1211), .A2(new_n749), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1122), .B2(new_n1013), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1118), .B(new_n1124), .C1(new_n1198), .C2(new_n1122), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n1015), .ZN(G381));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1207), .A2(new_n1233), .A3(new_n1209), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1037), .A2(new_n1013), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(new_n1009), .A3(new_n1012), .A4(new_n1010), .ZN(new_n1237));
  INV_X1    g1037(.A(G390), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n977), .A3(new_n1238), .ZN(new_n1239));
  OR3_X1    g1039(.A1(new_n1234), .A2(new_n1235), .A3(new_n1239), .ZN(G407));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(G343), .C2(new_n1234), .ZN(G409));
  NAND2_X1  g1041(.A1(new_n1206), .A2(G378), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n692), .A2(G213), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1231), .B2(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n709), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1230), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n858), .A3(new_n830), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(G384), .A3(new_n1230), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1199), .A2(new_n1014), .A3(new_n1196), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT124), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(KEYINPUT124), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1233), .B(new_n1197), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1251), .A4(new_n1255), .ZN(new_n1256));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  AND3_X1   g1057(.A1(new_n1237), .A2(new_n977), .A3(new_n1238), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1238), .B1(new_n1237), .B2(new_n977), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G387), .A2(G390), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1257), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1239), .A3(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1256), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1251), .A2(new_n1255), .A3(new_n1243), .A4(new_n1242), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1244), .A2(new_n1255), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n692), .A2(G213), .A3(G2897), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1249), .A2(new_n1250), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1269), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1265), .B(new_n1266), .C1(new_n1268), .C2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1244), .A2(new_n1279), .A3(new_n1251), .A4(new_n1255), .ZN(new_n1280));
  XOR2_X1   g1080(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1281));
  NAND4_X1  g1081(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1260), .A2(new_n1263), .A3(KEYINPUT126), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT126), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1276), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(new_n1234), .A2(new_n1242), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1251), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1234), .A2(new_n1251), .A3(new_n1242), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1285), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1285), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1290), .A2(new_n1285), .A3(new_n1297), .A4(new_n1291), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1293), .A2(new_n1296), .A3(new_n1298), .ZN(G402));
endmodule


