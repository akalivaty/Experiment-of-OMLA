//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT76), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(G211gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(G211gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT75), .B(G211gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT22), .B1(new_n212), .B2(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(G204gat), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(G197gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G204gat), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n211), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n226));
  OAI21_X1  g025(.A(G218gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n229), .A2(new_n210), .A3(new_n222), .A4(new_n217), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT3), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n237), .B2(KEYINPUT2), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G141gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G141gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n245), .A2(new_n247), .A3(G148gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n244), .B2(G148gat), .ZN(new_n250));
  INV_X1    g049(.A(G148gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT81), .B1(new_n251), .B2(G141gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(new_n247), .A3(G148gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n243), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n244), .A2(G148gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n251), .A2(G141gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n236), .A2(KEYINPUT79), .A3(new_n237), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n205), .B1(new_n233), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n243), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n269), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n231), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n231), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n261), .A2(KEYINPUT3), .A3(new_n270), .ZN(new_n283));
  INV_X1    g082(.A(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n269), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n224), .B2(new_n230), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(KEYINPUT3), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n285), .A2(KEYINPUT87), .A3(new_n205), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G22gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n229), .A2(new_n222), .A3(new_n217), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n284), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n293), .B2(new_n292), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n271), .B1(new_n295), .B2(new_n277), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n280), .A2(new_n296), .B1(new_n203), .B2(new_n204), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G78gat), .B(G106gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT86), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G50gat), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n291), .B1(new_n290), .B2(new_n297), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n304), .A2(KEYINPUT90), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT90), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT88), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n290), .A2(KEYINPUT88), .A3(new_n291), .A4(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n297), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G22gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315));
  INV_X1    g114(.A(new_n303), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n308), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT27), .B(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(new_n326), .B1(G183gat), .B2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT26), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT26), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n322), .A2(new_n336), .A3(new_n323), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n333), .B1(new_n330), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT23), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n330), .A2(KEYINPUT66), .A3(new_n339), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n346), .A2(KEYINPUT64), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OR3_X1    g149(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(KEYINPUT64), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n347), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT25), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n346), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(new_n349), .C1(G183gat), .C2(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(new_n343), .ZN(new_n357));
  INV_X1    g156(.A(new_n340), .ZN(new_n358));
  AND4_X1   g157(.A1(KEYINPUT25), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n338), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n360), .B2(new_n279), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n282), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n345), .A2(new_n353), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT25), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n368), .B2(new_n338), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n231), .B(new_n362), .C1(new_n369), .C2(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  OAI21_X1  g174(.A(KEYINPUT78), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377));
  INV_X1    g176(.A(new_n375), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n370), .A3(new_n375), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G127gat), .B(G134gat), .Z(new_n384));
  OR2_X1    g183(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G113gat), .B(G120gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n384), .B(new_n385), .C1(KEYINPUT1), .C2(new_n387), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT84), .B1(new_n271), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NOR4_X1   g193(.A1(new_n261), .A2(new_n391), .A3(new_n270), .A4(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT4), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n261), .B2(new_n270), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n278), .A2(new_n397), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  INV_X1    g203(.A(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(new_n395), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n271), .A2(new_n392), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n399), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT4), .B1(new_n393), .B2(new_n395), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n286), .B2(new_n391), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n398), .A2(new_n404), .A3(new_n399), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n403), .A2(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT0), .ZN(new_n419));
  XOR2_X1   g218(.A(G57gat), .B(G85gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT6), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n421), .B2(new_n417), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n417), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT6), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n383), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n308), .B(KEYINPUT91), .C1(new_n317), .C2(new_n318), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n321), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n416), .A2(new_n412), .A3(new_n414), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n393), .A2(new_n407), .A3(new_n395), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT5), .B1(new_n431), .B2(new_n399), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n432), .B2(new_n402), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n421), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT92), .B(new_n430), .C1(new_n432), .C2(new_n402), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n437), .A2(new_n422), .B1(KEYINPUT6), .B2(new_n424), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n378), .B1(new_n371), .B2(KEYINPUT37), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n231), .B1(new_n363), .B2(new_n364), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n282), .B(new_n362), .C1(new_n369), .C2(new_n361), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT37), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT38), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n381), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n365), .B2(new_n370), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT38), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(KEYINPUT93), .B(KEYINPUT38), .C1(new_n439), .C2(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n412), .A2(new_n398), .A3(new_n414), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n410), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n431), .B2(new_n399), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n455), .A3(new_n410), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n421), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n460), .A2(KEYINPUT40), .B1(new_n380), .B2(new_n382), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT40), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n435), .A2(new_n436), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n438), .A2(new_n452), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n392), .B1(new_n368), .B2(new_n338), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n392), .B(new_n338), .C1(new_n354), .C2(new_n359), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n469), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT32), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n360), .A2(new_n391), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n468), .B1(new_n478), .B2(new_n471), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT71), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n473), .B(KEYINPUT32), .C1(new_n474), .C2(new_n467), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT72), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n468), .A3(new_n471), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT34), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n484), .A2(new_n489), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n482), .A2(new_n488), .A3(new_n483), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT36), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n492), .A2(KEYINPUT36), .B1(new_n495), .B2(KEYINPUT73), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n464), .A2(new_n319), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n319), .A2(new_n426), .A3(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  INV_X1    g299(.A(new_n438), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n493), .A2(new_n494), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n502), .A2(new_n383), .A3(KEYINPUT35), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n319), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n429), .A2(new_n498), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT14), .B(G29gat), .Z(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G36gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  OR2_X1    g309(.A1(G43gat), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G43gat), .A2(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(G50gat), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n510), .B(new_n512), .C1(new_n515), .C2(G43gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT95), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n523), .A2(KEYINPUT95), .A3(G1gat), .ZN(new_n526));
  OAI221_X1 g325(.A(new_n521), .B1(G1gat), .B2(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT17), .B1(new_n514), .B2(new_n517), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n520), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n527), .B(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n518), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n533), .B(new_n518), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n532), .B(KEYINPUT13), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .A4(new_n534), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G197gat), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT11), .B(G169gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n537), .A2(new_n540), .A3(new_n547), .A4(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n505), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n423), .A2(new_n425), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g356(.A(G71gat), .ZN(new_n558));
  INV_X1    g357(.A(G78gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G127gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n562), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n561), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n533), .B1(KEYINPUT21), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n569), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n234), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n569), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n569), .A2(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT7), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n586), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n589), .B2(new_n593), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n518), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n520), .A2(new_n530), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n597), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT99), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605));
  INV_X1    g404(.A(new_n603), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n599), .B(new_n606), .C1(new_n600), .C2(new_n597), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n601), .A2(new_n605), .A3(new_n603), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT97), .Z(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n607), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n583), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n204), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n563), .B1(new_n595), .B2(new_n596), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n589), .A2(new_n593), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n590), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n571), .A2(new_n623), .A3(new_n594), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n571), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n620), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n628), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n628), .B2(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n553), .A2(new_n555), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n505), .A2(new_n552), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n383), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(G8gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT101), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT102), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n650), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n648), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(G1325gat));
  INV_X1    g457(.A(new_n643), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n496), .A2(new_n497), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n502), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n659), .B2(new_n662), .ZN(G1326gat));
  AND2_X1   g462(.A1(new_n321), .A2(new_n428), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n553), .A2(new_n664), .A3(new_n639), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR3_X1   g466(.A1(new_n583), .A2(new_n617), .A3(new_n638), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n553), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n506), .A3(new_n555), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT44), .B1(new_n505), .B2(new_n617), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n498), .A2(new_n429), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n500), .A2(new_n504), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n616), .A2(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n614), .A2(new_n678), .A3(new_n615), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n579), .A2(KEYINPUT103), .A3(new_n582), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT103), .B1(new_n579), .B2(new_n582), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(new_n552), .A3(new_n638), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n554), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n691), .ZN(G1328gat));
  INV_X1    g491(.A(new_n690), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(KEYINPUT105), .A3(new_n383), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  INV_X1    g494(.A(new_n383), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n690), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(G36gat), .A3(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n669), .A2(G36gat), .A3(new_n696), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1329gat));
  OAI21_X1  g500(.A(G43gat), .B1(new_n690), .B2(new_n660), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n669), .A2(G43gat), .A3(new_n502), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT47), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n704), .B(new_n706), .ZN(G1330gat));
  INV_X1    g506(.A(new_n515), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n670), .A2(new_n664), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n664), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n515), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n319), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n708), .B1(new_n693), .B2(new_n714), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n711), .A2(KEYINPUT48), .B1(new_n713), .B2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n638), .ZN(new_n717));
  NOR4_X1   g516(.A1(new_n505), .A2(new_n551), .A3(new_n618), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n555), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n383), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  INV_X1    g523(.A(new_n660), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n558), .B1(new_n718), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n502), .A2(G71gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n718), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n718), .A2(new_n664), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n583), .A2(new_n551), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n717), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n673), .B2(new_n683), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n554), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n676), .A2(new_n616), .A3(new_n732), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n676), .A2(KEYINPUT51), .A3(new_n616), .A4(new_n732), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT107), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n555), .A2(new_n584), .A3(new_n638), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(G1336gat));
  AOI21_X1  g545(.A(new_n585), .B1(new_n736), .B2(new_n383), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n717), .A2(G92gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n383), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n741), .B2(new_n742), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n676), .B2(new_n616), .ZN(new_n754));
  INV_X1    g553(.A(new_n682), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n505), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n383), .B(new_n734), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n752), .B1(new_n758), .B2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(new_n749), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n751), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n751), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(G1337gat));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n737), .B2(new_n660), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n736), .A2(KEYINPUT110), .A3(new_n725), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(G99gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n502), .A2(G99gat), .A3(new_n717), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT111), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n744), .B2(new_n772), .ZN(G1338gat));
  INV_X1    g572(.A(G106gat), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n736), .B2(new_n664), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n714), .A2(new_n774), .A3(new_n638), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(new_n743), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n774), .B1(new_n736), .B2(new_n714), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n743), .A2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n779), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n538), .A2(new_n539), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n532), .B1(new_n531), .B2(new_n534), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n546), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(new_n550), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n677), .A2(new_n679), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n628), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n626), .A2(new_n627), .A3(new_n620), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n628), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n793), .B2(new_n635), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n795), .B(new_n634), .C1(new_n628), .C2(new_n792), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT55), .B(new_n791), .C1(new_n794), .C2(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n636), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n799), .A2(new_n551), .A3(new_n636), .A4(new_n800), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n638), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(new_n804), .B1(new_n677), .B2(new_n679), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n687), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n639), .A2(new_n552), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n502), .B(new_n664), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n555), .A2(new_n696), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n552), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n554), .B1(new_n806), .B2(new_n807), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n319), .A2(new_n492), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n696), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT113), .Z(new_n817));
  INV_X1    g616(.A(G113gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n551), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n812), .B2(new_n717), .ZN(new_n821));
  INV_X1    g620(.A(G120gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n817), .A2(new_n822), .A3(new_n638), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1341gat));
  NAND3_X1  g623(.A1(new_n811), .A2(G127gat), .A3(new_n688), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(new_n583), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n568), .B1(new_n816), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(G1342gat));
  OAI21_X1  g629(.A(G134gat), .B1(new_n812), .B2(new_n617), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n815), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n832), .A2(G134gat), .A3(new_n383), .A4(new_n617), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT56), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1343gat));
  NOR2_X1   g634(.A1(new_n725), .A2(new_n809), .ZN(new_n836));
  XOR2_X1   g635(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n837));
  NAND2_X1  g636(.A1(new_n797), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(new_n551), .A3(new_n636), .A4(new_n800), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n804), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n839), .B2(new_n804), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n617), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n801), .B2(new_n788), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n827), .B1(new_n552), .B2(new_n639), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n664), .A2(KEYINPUT57), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n806), .A2(new_n807), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n714), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n846), .A2(new_n847), .B1(new_n849), .B2(KEYINPUT115), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n551), .B(new_n836), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n245), .A2(new_n247), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n725), .A2(new_n319), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n814), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n696), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(G141gat), .A3(new_n552), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n852), .A2(new_n862), .A3(new_n853), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n852), .B2(new_n853), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(new_n859), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(G1344gat));
  INV_X1    g666(.A(new_n858), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n251), .A3(new_n638), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n836), .B1(new_n850), .B2(new_n851), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n717), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(KEYINPUT59), .A3(new_n251), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n839), .A2(new_n804), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n616), .B1(new_n875), .B2(new_n841), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n616), .A2(new_n787), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n801), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n827), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n807), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n664), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n848), .A2(new_n714), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT57), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n638), .A3(new_n836), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n869), .B1(new_n872), .B2(new_n886), .ZN(G1345gat));
  OAI21_X1  g686(.A(G155gat), .B1(new_n870), .B2(new_n687), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n234), .A3(new_n583), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n870), .B2(new_n681), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n857), .A2(new_n235), .A3(new_n696), .A4(new_n616), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n555), .A2(new_n696), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n808), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n552), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT121), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n555), .B1(new_n806), .B2(new_n807), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n383), .A3(new_n815), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n328), .A3(new_n551), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(G1348gat));
  OAI21_X1  g703(.A(G176gat), .B1(new_n897), .B2(new_n717), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n329), .A3(new_n638), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT122), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n808), .A2(new_n688), .A3(new_n896), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n583), .A2(new_n322), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n909), .A2(G183gat), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n911), .B(new_n912), .Z(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n897), .B2(new_n617), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n323), .A3(new_n680), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(G1351gat));
  AND3_X1   g719(.A1(new_n855), .A2(new_n900), .A3(new_n383), .ZN(new_n921));
  AOI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n551), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n660), .A2(new_n896), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n882), .A2(new_n884), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n552), .A2(new_n219), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n214), .A3(new_n638), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT62), .Z(new_n929));
  OAI21_X1  g728(.A(G204gat), .B1(new_n924), .B2(new_n717), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT125), .ZN(G1353gat));
  INV_X1    g731(.A(new_n212), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n921), .A2(new_n933), .A3(new_n583), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n882), .A2(new_n583), .A3(new_n884), .A4(new_n923), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(G1354gat));
  NAND3_X1  g739(.A1(new_n921), .A2(new_n207), .A3(new_n680), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n942), .A2(new_n943), .A3(new_n617), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n944), .B2(new_n207), .ZN(G1355gat));
endmodule


