//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n220), .A2(new_n207), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT0), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n226), .B1(new_n225), .B2(new_n224), .C1(new_n216), .C2(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n218), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  AND2_X1   g0044(.A1(G1), .A2(G13), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n245), .B1(new_n208), .B2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT70), .A2(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT8), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(new_n207), .A3(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n246), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n206), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n256), .A2(new_n258), .B1(G50), .B2(new_n255), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(G226), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(G222), .B1(G77), .B2(new_n271), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G1698), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT67), .B(G223), .Z(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n273), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(KEYINPUT69), .A3(new_n221), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n245), .B2(new_n264), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n280), .B2(new_n281), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n268), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(G169), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n261), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT71), .B(new_n261), .C1(new_n291), .C2(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G68), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n254), .A2(G20), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(KEYINPUT78), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(KEYINPUT78), .ZN(new_n304));
  INV_X1    g0104(.A(new_n256), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n299), .B1(new_n206), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n246), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n299), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n207), .A2(G33), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT77), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n307), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n276), .A2(G226), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n320), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n288), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n263), .B1(new_n267), .B2(G238), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n319), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n319), .A3(new_n328), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n331), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n318), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT79), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(new_n331), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n340), .B(new_n344), .C1(new_n341), .C2(new_n329), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(G179), .A3(new_n331), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n337), .B1(new_n347), .B2(new_n318), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n257), .A2(G77), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n256), .A2(new_n349), .B1(G77), .B2(new_n255), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(new_n311), .B1(new_n207), .B2(new_n310), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  INV_X1    g0153(.A(new_n250), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n308), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n263), .B1(new_n267), .B2(G244), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n276), .A2(G232), .A3(new_n321), .ZN(new_n362));
  INV_X1    g0162(.A(G107), .ZN(new_n363));
  INV_X1    g0163(.A(G238), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n362), .B1(new_n363), .B2(new_n276), .C1(new_n277), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n365), .B2(new_n288), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n366), .A2(new_n335), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(G200), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n359), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(G179), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n338), .B2(new_n366), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(new_n358), .ZN(new_n372));
  INV_X1    g0172(.A(new_n350), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n298), .A2(new_n348), .A3(new_n369), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n290), .A2(G200), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT9), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT73), .B1(new_n261), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n261), .A2(new_n378), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(G190), .B(new_n268), .C1(new_n283), .C2(new_n289), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n261), .A2(KEYINPUT73), .A3(new_n378), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n377), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT10), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT74), .B1(new_n384), .B2(KEYINPUT10), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(KEYINPUT74), .A3(KEYINPUT10), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(G223), .B(new_n321), .C1(new_n269), .C2(new_n270), .ZN(new_n390));
  OAI211_X1 g0190(.A(G226), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n288), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n262), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT82), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n393), .B2(new_n288), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT82), .ZN(new_n402));
  AOI21_X1  g0202(.A(G169), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(G179), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT83), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n271), .B2(new_n207), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n269), .A2(new_n270), .A3(new_n407), .A4(G20), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G58), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n299), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n411), .B2(new_n201), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n250), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n246), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n274), .A2(new_n207), .A3(new_n275), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n407), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n275), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n414), .B1(new_n422), .B2(G68), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT80), .B1(new_n423), .B2(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n299), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT80), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n425), .A2(new_n426), .A3(new_n414), .A4(new_n417), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n418), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n248), .A2(new_n257), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n429), .A2(new_n256), .B1(new_n255), .B2(new_n248), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT81), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n399), .B(new_n396), .C1(new_n288), .C2(new_n393), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT82), .B1(new_n394), .B2(new_n397), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n338), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT83), .ZN(new_n437));
  INV_X1    g0237(.A(new_n404), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n405), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT18), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n405), .A2(new_n433), .A3(new_n442), .A4(new_n439), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n333), .B1(new_n434), .B2(new_n435), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n401), .A2(new_n335), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n428), .A3(new_n432), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n446), .A2(KEYINPUT17), .A3(new_n428), .A4(new_n432), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n441), .A2(new_n443), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n376), .A2(new_n389), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n206), .A2(G33), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n246), .A2(new_n255), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G107), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n207), .A2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n254), .A2(new_n457), .A3(KEYINPUT25), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT25), .B1(new_n254), .B2(new_n457), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT93), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n460), .B2(new_n458), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n207), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n276), .A2(new_n465), .A3(new_n207), .A4(G87), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n363), .A2(KEYINPUT23), .A3(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT23), .B1(new_n363), .B2(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n468), .A2(new_n469), .B1(G20), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(KEYINPUT24), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n308), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT24), .B1(new_n467), .B2(new_n472), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n456), .B(new_n462), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n321), .C1(new_n269), .C2(new_n270), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT94), .A3(new_n288), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(new_n485), .B1(new_n245), .B2(new_n264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n206), .A2(G45), .ZN(new_n487));
  OR2_X1    g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NAND2_X1  g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n486), .A2(G264), .B1(G274), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT94), .B1(new_n481), .B2(new_n288), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT95), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n493), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT95), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n482), .A4(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n481), .A2(new_n288), .B1(new_n486), .B2(G264), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n490), .A2(G274), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n292), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n477), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n497), .A3(new_n335), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n333), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n477), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT96), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(KEYINPUT96), .A3(new_n477), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n454), .A2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n255), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G20), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(G33), .ZN(new_n519));
  INV_X1    g0319(.A(G283), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(KEYINPUT85), .A2(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT85), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n518), .B1(new_n525), .B2(G20), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT20), .B1(new_n526), .B2(new_n308), .ZN(new_n527));
  AND2_X1   g0327(.A1(KEYINPUT85), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(KEYINPUT85), .A2(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n521), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n518), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT20), .B(new_n308), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n517), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT91), .B(G303), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n271), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n321), .C1(new_n269), .C2(new_n270), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT92), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n538), .A2(KEYINPUT92), .A3(new_n539), .A4(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n288), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n486), .A2(G270), .B1(G274), .B2(new_n490), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n536), .A2(G169), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n547), .A2(new_n292), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n536), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n536), .A2(KEYINPUT21), .A3(G169), .A4(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(new_n536), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n547), .A2(G190), .ZN(new_n554));
  AOI21_X1  g0354(.A(G200), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n284), .A2(new_n221), .ZN(new_n558));
  OAI21_X1  g0358(.A(G250), .B1(new_n484), .B2(G1), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT88), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT88), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n265), .A2(new_n561), .A3(G250), .A4(new_n487), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n560), .A2(new_n562), .B1(G274), .B2(new_n485), .ZN(new_n563));
  OAI211_X1 g0363(.A(G238), .B(new_n321), .C1(new_n269), .C2(new_n270), .ZN(new_n564));
  OAI211_X1 g0364(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n470), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n288), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n567), .A3(G190), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT90), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT90), .A4(G190), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n207), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n311), .B1(new_n522), .B2(new_n523), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(KEYINPUT19), .ZN(new_n575));
  NAND3_X1  g0375(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n576), .A2(new_n207), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n528), .A2(new_n529), .A3(G107), .ZN(new_n578));
  XNOR2_X1  g0378(.A(KEYINPUT89), .B(G87), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n308), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n255), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n351), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n246), .A2(G87), .A3(new_n255), .A4(new_n453), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n333), .B1(new_n563), .B2(new_n567), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n563), .A2(new_n567), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n563), .A2(new_n567), .A3(G179), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n581), .B(new_n583), .C1(new_n351), .C2(new_n454), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n572), .A2(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n582), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n454), .B2(new_n594), .ZN(new_n596));
  OR2_X1    g0396(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n597));
  NAND2_X1  g0397(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n598));
  AND2_X1   g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  NOR2_X1   g0399(.A1(G97), .A2(G107), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n528), .A2(new_n529), .ZN(new_n602));
  AND2_X1   g0402(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n603));
  NOR2_X1   g0403(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n363), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G20), .ZN(new_n607));
  OAI21_X1  g0407(.A(G107), .B1(new_n406), .B2(new_n408), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n250), .A2(G77), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n596), .B1(new_n610), .B2(new_n308), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT4), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G1698), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(G244), .C1(new_n270), .C2(new_n269), .ZN(new_n615));
  INV_X1    g0415(.A(G244), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n274), .B2(new_n275), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n531), .C1(new_n617), .C2(KEYINPUT4), .ZN(new_n618));
  OAI21_X1  g0418(.A(G250), .B1(new_n269), .B2(new_n270), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n321), .B1(new_n619), .B2(KEYINPUT4), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n288), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n489), .ZN(new_n622));
  NOR2_X1   g0422(.A1(KEYINPUT5), .A2(G41), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n485), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(G257), .A3(new_n265), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n501), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G169), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(KEYINPUT86), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n625), .A2(new_n501), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n621), .A2(new_n630), .A3(new_n292), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n612), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n621), .A2(new_n630), .A3(new_n632), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT87), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n621), .A2(new_n630), .A3(new_n637), .A4(new_n632), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n333), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n621), .A2(new_n627), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n611), .B1(new_n335), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n593), .B(new_n634), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n557), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n452), .A2(new_n513), .A3(new_n643), .ZN(G372));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(new_n633), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n646), .A2(new_n611), .A3(new_n628), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n593), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n591), .A2(new_n592), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n593), .B2(new_n647), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT96), .B1(new_n508), .B2(new_n477), .ZN(new_n653));
  AOI211_X1 g0453(.A(new_n510), .B(new_n476), .C1(new_n506), .C2(new_n507), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n548), .A2(new_n549), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n550), .A2(new_n536), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n552), .A3(new_n656), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n653), .A2(new_n654), .B1(new_n657), .B2(new_n505), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n658), .B2(new_n642), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n452), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n345), .A2(new_n346), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n344), .B1(new_n332), .B2(new_n340), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n318), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n663), .A2(new_n375), .ZN(new_n664));
  INV_X1    g0464(.A(new_n337), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n449), .A3(new_n450), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n441), .B(new_n443), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n388), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n668), .A2(new_n386), .B1(KEYINPUT10), .B2(new_n384), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(new_n669), .B1(new_n296), .B2(new_n297), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n660), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT97), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  OAI21_X1  g0474(.A(G213), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n676), .A3(new_n674), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT97), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n672), .B(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT98), .B1(new_n679), .B2(KEYINPUT27), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n675), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n553), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT99), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n557), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n684), .B2(new_n557), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n657), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  AOI211_X1 g0489(.A(new_n689), .B(new_n675), .C1(new_n677), .C2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n476), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n513), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n338), .B1(new_n494), .B2(new_n497), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n476), .B1(new_n693), .B2(new_n503), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n694), .B2(new_n682), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n688), .A2(new_n695), .A3(G330), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n505), .A2(new_n682), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n657), .A2(new_n682), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n513), .A2(new_n691), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(G399));
  NAND3_X1  g0501(.A1(new_n578), .A2(new_n515), .A3(new_n579), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  INV_X1    g0503(.A(new_n223), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n703), .A2(new_n206), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n220), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND2_X1  g0509(.A1(new_n572), .A2(new_n587), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n634), .B(new_n710), .C1(new_n639), .C2(new_n641), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n551), .A2(new_n694), .A3(new_n552), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n712), .B(new_n713), .C1(new_n653), .C2(new_n654), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n690), .B1(new_n714), .B2(new_n652), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT103), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n659), .A2(new_n682), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(KEYINPUT103), .B(KEYINPUT29), .C1(new_n659), .C2(new_n682), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n513), .A2(new_n643), .A3(new_n682), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(new_n588), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n500), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT101), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT102), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n640), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n500), .A3(KEYINPUT101), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n550), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n729), .B2(new_n730), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n729), .A2(new_n730), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n550), .A3(new_n728), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n725), .A2(G179), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n502), .A3(new_n635), .A4(new_n547), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n724), .B1(new_n740), .B2(new_n690), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n724), .A3(new_n690), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n722), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n709), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n253), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n705), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n688), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(G330), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n686), .A2(new_n754), .A3(new_n687), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT107), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n688), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n704), .A2(new_n271), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n515), .B2(new_n704), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n707), .A2(G45), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n243), .B2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n704), .A2(new_n276), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n763), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n221), .B1(G20), .B2(new_n338), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n207), .A2(G190), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n207), .A2(new_n335), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n292), .A2(new_n333), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n292), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n202), .B1(new_n784), .B2(new_n310), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n207), .B1(new_n775), .B2(G190), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n781), .A2(new_n772), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n276), .B1(new_n786), .B2(new_n594), .C1(new_n299), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n780), .A2(new_n783), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n785), .B(new_n788), .C1(G58), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n292), .A2(G200), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT105), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n780), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(new_n579), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n773), .A3(new_n774), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G107), .ZN(new_n798));
  AND4_X1   g0598(.A1(new_n779), .A2(new_n791), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n776), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n797), .A2(G283), .B1(G329), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT106), .Z(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n271), .B1(new_n786), .B2(new_n803), .C1(new_n782), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n787), .ZN(new_n806));
  NOR2_X1   g0606(.A1(KEYINPUT33), .A2(G317), .ZN(new_n807));
  AND2_X1   g0607(.A1(KEYINPUT33), .A2(G317), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n784), .C1(new_n811), .C2(new_n789), .ZN(new_n812));
  INV_X1    g0612(.A(new_n794), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n805), .B(new_n812), .C1(G303), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n799), .B1(new_n802), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n769), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n771), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n761), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n756), .B1(new_n752), .B2(new_n818), .ZN(G396));
  INV_X1    g0619(.A(new_n745), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT109), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n374), .A2(new_n690), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT109), .B1(new_n359), .B2(new_n682), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n369), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n375), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n371), .A2(new_n374), .A3(new_n682), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n718), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n752), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n820), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n752), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n769), .A2(new_n757), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n310), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n797), .A2(G87), .B1(G311), .B2(new_n800), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n363), .B2(new_n794), .ZN(new_n836));
  INV_X1    g0636(.A(new_n784), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G283), .A2(new_n806), .B1(new_n837), .B2(G116), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n803), .B2(new_n789), .ZN(new_n839));
  INV_X1    g0639(.A(G303), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n271), .B1(new_n786), .B2(new_n594), .C1(new_n782), .C2(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G143), .A2(new_n790), .B1(new_n806), .B2(G150), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n844), .B2(new_n782), .C1(new_n777), .C2(new_n784), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n276), .B1(new_n410), .B2(new_n786), .C1(new_n776), .C2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n797), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n202), .B2(new_n794), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT108), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n842), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n834), .B1(new_n816), .B2(new_n855), .C1(new_n828), .C2(new_n758), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n831), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR3_X1   g0658(.A1(new_n221), .A2(new_n207), .A3(new_n515), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n606), .B2(KEYINPUT35), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(KEYINPUT35), .B2(new_n606), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT36), .ZN(new_n862));
  OR3_X1    g0662(.A1(new_n220), .A2(new_n310), .A3(new_n411), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n202), .A2(G68), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n206), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n681), .ZN(new_n867));
  INV_X1    g0667(.A(new_n430), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n428), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n451), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n433), .A2(new_n681), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n440), .A2(new_n871), .A3(new_n447), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n447), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n428), .A2(new_n868), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n870), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n318), .A2(new_n690), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n665), .A2(new_n663), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n318), .B(new_n690), .C1(new_n347), .C2(new_n337), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n827), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n887), .A2(new_n742), .A3(new_n743), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT111), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n742), .A3(new_n743), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT111), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n883), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n870), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(new_n872), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n440), .A2(new_n447), .A3(new_n872), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n451), .A2(new_n896), .B1(new_n898), .B2(new_n873), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n895), .B1(KEYINPUT38), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n889), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n452), .A2(new_n744), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n754), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n347), .A2(new_n318), .A3(new_n682), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n895), .B(new_n908), .C1(KEYINPUT38), .C2(new_n899), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n870), .A2(new_n880), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n913), .B2(new_n895), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT110), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n441), .A2(new_n443), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n867), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n885), .A2(new_n886), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n920));
  INV_X1    g0720(.A(new_n593), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n713), .C1(new_n653), .C2(new_n654), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n690), .B(new_n827), .C1(new_n923), .C2(new_n652), .ZN(new_n924));
  INV_X1    g0724(.A(new_n826), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n916), .B(new_n918), .C1(new_n926), .C2(new_n883), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n919), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n659), .A2(new_n682), .A3(new_n828), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n826), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n913), .A2(new_n895), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n916), .B1(new_n933), .B2(new_n918), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n452), .B(new_n716), .C1(new_n720), .C2(new_n721), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n670), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n905), .A2(new_n938), .B1(new_n206), .B2(new_n749), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n905), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n866), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n690), .A2(new_n585), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT112), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n593), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n649), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n697), .B1(new_n700), .B2(KEYINPUT42), .ZN(new_n947));
  INV_X1    g0747(.A(new_n920), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n612), .A2(new_n690), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT42), .B1(new_n700), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n634), .B2(new_n690), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n946), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n696), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n952), .B1(new_n634), .B2(new_n682), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n959), .B(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n705), .B(KEYINPUT41), .Z(new_n965));
  NAND3_X1  g0765(.A1(new_n700), .A2(new_n697), .A3(new_n961), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT45), .Z(new_n967));
  AOI21_X1  g0767(.A(new_n961), .B1(new_n700), .B2(new_n697), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n960), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n967), .A2(new_n696), .A3(new_n970), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n700), .B1(new_n695), .B2(new_n699), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n753), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n746), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n965), .B1(new_n978), .B2(new_n747), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n964), .B1(new_n979), .B2(new_n751), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n767), .A2(new_n235), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n770), .B1(new_n223), .B2(new_n351), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n752), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n276), .B1(new_n784), .B2(new_n202), .ZN(new_n984));
  INV_X1    g0784(.A(new_n782), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G143), .A2(new_n985), .B1(new_n790), .B2(G150), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n777), .B2(new_n787), .ZN(new_n987));
  INV_X1    g0787(.A(new_n786), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n984), .B(new_n987), .C1(G68), .C2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n794), .A2(new_n410), .B1(new_n776), .B2(new_n844), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G77), .B2(new_n797), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n794), .A2(new_n515), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n796), .A2(new_n602), .B1(new_n995), .B2(new_n776), .ZN(new_n996));
  INV_X1    g0796(.A(new_n537), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n789), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n787), .A2(new_n803), .B1(new_n784), .B2(new_n520), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT114), .B(G311), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n271), .B1(new_n786), .B2(new_n363), .C1(new_n782), .C2(new_n1000), .ZN(new_n1001));
  NOR4_X1   g0801(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n989), .A2(new_n991), .B1(new_n994), .B2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT47), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n816), .B1(new_n1003), .B2(KEYINPUT47), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n983), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n945), .B2(new_n760), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n980), .A2(new_n1007), .ZN(G387));
  INV_X1    g0808(.A(new_n977), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n746), .A2(new_n976), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n705), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n695), .A2(new_n760), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n353), .A2(G50), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT50), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n484), .B1(new_n299), .B2(new_n310), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n703), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n766), .B1(new_n232), .B2(new_n484), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n703), .A2(new_n762), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n223), .A2(G107), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n770), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n782), .A2(new_n777), .B1(new_n784), .B2(new_n299), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n271), .B(new_n1022), .C1(G50), .C2(new_n790), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n813), .A2(G77), .B1(new_n800), .B2(G150), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n351), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n248), .A2(new_n806), .B1(new_n988), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n797), .A2(G97), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n794), .A2(new_n803), .B1(new_n520), .B2(new_n786), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n997), .A2(new_n784), .B1(new_n782), .B2(new_n811), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1000), .A2(new_n787), .B1(new_n789), .B2(new_n995), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(KEYINPUT48), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(KEYINPUT48), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n276), .B1(new_n797), .B2(G116), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n804), .C2(new_n776), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1028), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n832), .B1(new_n1039), .B2(new_n769), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1021), .A2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1011), .B1(new_n750), .B2(new_n976), .C1(new_n1012), .C2(new_n1041), .ZN(G393));
  OAI221_X1 g0842(.A(new_n770), .B1(new_n223), .B2(new_n602), .C1(new_n240), .C2(new_n767), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT115), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n832), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n782), .A2(new_n995), .B1(new_n789), .B2(new_n810), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT52), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1047), .A2(new_n1048), .B1(new_n776), .B2(new_n811), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G283), .B2(new_n813), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n784), .A2(new_n803), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n271), .B1(new_n997), .B2(new_n787), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G116), .C2(new_n988), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n798), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n797), .A2(G87), .B1(G143), .B2(new_n800), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n276), .B1(new_n784), .B2(new_n353), .C1(new_n202), .C2(new_n787), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G77), .B2(new_n988), .ZN(new_n1058));
  INV_X1    g0858(.A(G150), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n782), .A2(new_n1059), .B1(new_n789), .B2(new_n777), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n813), .A2(G68), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1056), .A2(new_n1058), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n816), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1046), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n759), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n961), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n974), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n750), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n705), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n974), .B2(new_n977), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1009), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G390));
  OAI21_X1  g0874(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n909), .C1(new_n931), .C2(new_n907), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n925), .B1(new_n715), .B2(new_n825), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n900), .B(new_n906), .C1(new_n1077), .C2(new_n929), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n887), .A2(new_n742), .A3(G330), .A4(new_n743), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(KEYINPUT116), .B(new_n1079), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1075), .A2(new_n909), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n930), .A2(new_n826), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n907), .B1(new_n1084), .B2(new_n919), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1078), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1079), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1080), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1075), .A2(new_n757), .A3(new_n909), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n833), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n752), .B1(new_n248), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n276), .B1(new_n813), .B2(G87), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT117), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n789), .A2(new_n515), .B1(new_n784), .B2(new_n602), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n782), .A2(new_n520), .B1(new_n787), .B2(new_n363), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G77), .C2(new_n988), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(new_n852), .C1(new_n803), .C2(new_n776), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G132), .A2(new_n790), .B1(new_n837), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n844), .B2(new_n787), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n796), .A2(new_n202), .B1(new_n1104), .B2(new_n776), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n276), .B1(new_n786), .B2(new_n777), .C1(new_n782), .C2(new_n1106), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n813), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1095), .A2(new_n1099), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1093), .B1(new_n1111), .B2(new_n769), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1090), .A2(new_n751), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n742), .A2(G330), .A3(new_n743), .A4(new_n828), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n929), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1077), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n1079), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n888), .A2(G330), .B1(new_n1114), .B2(new_n929), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n1084), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n452), .A2(new_n744), .A3(G330), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n936), .A2(new_n670), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1089), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1080), .B(new_n1122), .C1(new_n1081), .C2(new_n1088), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n705), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1113), .A2(new_n1126), .ZN(G378));
  NOR2_X1   g0927(.A1(new_n867), .A2(new_n260), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n294), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n389), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1128), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n669), .A2(new_n294), .A3(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n928), .B2(new_n934), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n918), .B1(new_n926), .B2(new_n883), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT110), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n1137), .A3(new_n927), .A4(new_n915), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(G330), .B1(new_n894), .B2(new_n901), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1139), .A2(new_n1144), .A3(new_n1142), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1121), .B(KEYINPUT122), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1146), .A2(new_n1147), .B1(new_n1125), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT123), .B1(new_n1149), .B2(KEYINPUT57), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1070), .B1(new_n1149), .B2(KEYINPUT57), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT123), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1139), .A2(new_n1144), .A3(new_n1142), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1144), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1152), .B(new_n1153), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1150), .A2(new_n1151), .A3(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n276), .A2(G41), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n789), .B2(new_n363), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n790), .A2(KEYINPUT118), .A3(G107), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(G77), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n797), .A2(G58), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n520), .C2(new_n776), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1160), .B1(new_n985), .B2(G116), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G97), .A2(new_n806), .B1(new_n837), .B2(new_n1025), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n299), .C2(new_n786), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1161), .B1(new_n1171), .B2(KEYINPUT58), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT119), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n797), .C2(G159), .ZN(new_n1174));
  INV_X1    g0974(.A(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n776), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n784), .A2(new_n844), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n782), .A2(new_n1104), .B1(new_n787), .B2(new_n849), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G150), .C2(new_n988), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n794), .A2(new_n1100), .B1(new_n1106), .B2(new_n789), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1184), .B2(KEYINPUT59), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1185), .A2(new_n1186), .B1(KEYINPUT58), .B2(new_n1171), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1173), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n769), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n752), .B1(G50), .B2(new_n1092), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1137), .B2(new_n757), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n751), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1159), .A2(new_n1196), .ZN(G375));
  INV_X1    g0997(.A(new_n1119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n929), .A2(new_n757), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n752), .B1(G68), .B2(new_n1092), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n797), .A2(G77), .B1(G303), .B2(new_n800), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n594), .B2(new_n794), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G294), .A2(new_n985), .B1(new_n837), .B2(G107), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n988), .A2(new_n1025), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n790), .A2(G283), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n276), .B1(new_n806), .B2(G116), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n782), .A2(new_n849), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n813), .A2(G159), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n800), .A2(G128), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1166), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n806), .A2(new_n1101), .B1(new_n837), .B2(G150), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n271), .B1(new_n790), .B2(G137), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n202), .C2(new_n786), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1202), .A2(new_n1207), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1200), .B1(new_n1216), .B2(new_n769), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1198), .A2(new_n751), .B1(new_n1199), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n965), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1123), .A2(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT125), .ZN(G381));
  NAND2_X1  g1023(.A1(G378), .A2(KEYINPUT126), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1126), .A2(new_n1225), .A3(new_n1113), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G375), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1073), .A2(new_n980), .A3(new_n1007), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(G407));
  AND2_X1   g1032(.A1(new_n689), .A2(G213), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1228), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  NAND2_X1  g1035(.A1(G387), .A2(G390), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1229), .ZN(new_n1237));
  AND2_X1   g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1236), .A3(new_n1229), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n1121), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1246), .B(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1122), .A2(new_n1070), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(KEYINPUT60), .C2(new_n1221), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G384), .B1(new_n1250), .B2(new_n1218), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(G384), .A3(new_n1218), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1159), .A2(G378), .A3(new_n1196), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1149), .A2(new_n1219), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1196), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1224), .A2(new_n1257), .A3(new_n1226), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1233), .B(new_n1254), .C1(new_n1255), .C2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1245), .B1(new_n1259), .B2(KEYINPUT63), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1233), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1253), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G2897), .B(new_n1233), .C1(new_n1262), .C2(new_n1251), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1233), .A2(G2897), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1252), .A2(new_n1253), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT63), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1254), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1260), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1261), .A2(new_n1272), .A3(new_n1268), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1243), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1261), .B2(new_n1268), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1244), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1240), .B1(new_n1236), .B2(new_n1229), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1271), .B1(new_n1276), .B2(new_n1279), .ZN(G405));
  OAI21_X1  g1080(.A(new_n1254), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1242), .A2(new_n1268), .A3(new_n1244), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1255), .B1(new_n1284), .B2(new_n1227), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1283), .B(new_n1285), .Z(G402));
endmodule


