

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U324 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U325 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U326 ( .A(n457), .B(n326), .ZN(n523) );
  XNOR2_X1 U327 ( .A(n436), .B(n323), .ZN(n324) );
  AND2_X1 U328 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n348) );
  XNOR2_X1 U330 ( .A(n349), .B(n348), .ZN(n389) );
  XNOR2_X1 U331 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U332 ( .A(n378), .B(n299), .ZN(n303) );
  NOR2_X1 U333 ( .A1(n439), .A2(n473), .ZN(n440) );
  INV_X1 U334 ( .A(G106GAT), .ZN(n382) );
  XNOR2_X1 U335 ( .A(n359), .B(n292), .ZN(n323) );
  INV_X1 U336 ( .A(KEYINPUT64), .ZN(n422) );
  XNOR2_X1 U337 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U338 ( .A(KEYINPUT37), .B(KEYINPUT110), .ZN(n496) );
  XNOR2_X1 U339 ( .A(n423), .B(n422), .ZN(n568) );
  XNOR2_X1 U340 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U341 ( .A(n497), .B(n496), .ZN(n519) );
  XNOR2_X1 U342 ( .A(n499), .B(KEYINPUT38), .ZN(n507) );
  XNOR2_X1 U343 ( .A(n462), .B(G176GAT), .ZN(n463) );
  XNOR2_X1 U344 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U346 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n312) );
  XOR2_X1 U348 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n296) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n378) );
  NAND2_X1 U351 ( .A1(G230GAT), .A2(G233GAT), .ZN(n298) );
  INV_X1 U352 ( .A(KEYINPUT76), .ZN(n297) );
  XOR2_X1 U353 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n301) );
  XOR2_X1 U354 ( .A(G106GAT), .B(G78GAT), .Z(n424) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G64GAT), .Z(n318) );
  XNOR2_X1 U356 ( .A(n424), .B(n318), .ZN(n300) );
  XOR2_X1 U357 ( .A(n301), .B(n300), .Z(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n310) );
  XNOR2_X1 U359 ( .A(G120GAT), .B(G148GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n304), .B(G57GAT), .ZN(n409) );
  XOR2_X1 U361 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n306) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(KEYINPUT75), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n355) );
  XNOR2_X1 U364 ( .A(n409), .B(n355), .ZN(n308) );
  XNOR2_X1 U365 ( .A(G204GAT), .B(G92GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n393) );
  XNOR2_X1 U367 ( .A(KEYINPUT41), .B(n393), .ZN(n548) );
  XOR2_X1 U368 ( .A(KEYINPUT19), .B(KEYINPUT92), .Z(n314) );
  XNOR2_X1 U369 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(G169GAT), .B(n315), .Z(n457) );
  XOR2_X1 U372 ( .A(G92GAT), .B(KEYINPUT87), .Z(n317) );
  XNOR2_X1 U373 ( .A(G36GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n368) );
  XNOR2_X1 U375 ( .A(n368), .B(n318), .ZN(n325) );
  XNOR2_X1 U376 ( .A(G211GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n319), .B(KEYINPUT21), .ZN(n320) );
  XOR2_X1 U378 ( .A(n320), .B(KEYINPUT95), .Z(n322) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n436) );
  XOR2_X1 U381 ( .A(G8GAT), .B(G183GAT), .Z(n359) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n327), .B(KEYINPUT7), .ZN(n381) );
  XOR2_X1 U385 ( .A(n381), .B(KEYINPUT71), .Z(n329) );
  NAND2_X1 U386 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT73), .Z(n331) );
  XNOR2_X1 U389 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U392 ( .A(G1GAT), .B(G141GAT), .Z(n335) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(G197GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G50GAT), .Z(n340) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(G22GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n338), .B(KEYINPUT72), .ZN(n356) );
  XNOR2_X1 U399 ( .A(G113GAT), .B(n356), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U401 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U402 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n345), .B(G36GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n557) );
  NOR2_X1 U407 ( .A1(n557), .A2(n548), .ZN(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n351) );
  XNOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n367) );
  XOR2_X1 U411 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n353) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(n354), .B(KEYINPUT90), .Z(n358) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U417 ( .A(G1GAT), .B(G127GAT), .Z(n417) );
  XOR2_X1 U418 ( .A(n359), .B(n417), .Z(n361) );
  XNOR2_X1 U419 ( .A(G155GAT), .B(G57GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U421 ( .A(n363), .B(n362), .Z(n365) );
  XNOR2_X1 U422 ( .A(G211GAT), .B(G78GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U424 ( .A(n367), .B(n366), .Z(n576) );
  XOR2_X1 U425 ( .A(G50GAT), .B(KEYINPUT82), .Z(n425) );
  XOR2_X1 U426 ( .A(n368), .B(n425), .Z(n370) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n387) );
  XOR2_X1 U429 ( .A(KEYINPUT84), .B(KEYINPUT66), .Z(n372) );
  XNOR2_X1 U430 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT10), .B(KEYINPUT83), .Z(n374) );
  XNOR2_X1 U433 ( .A(KEYINPUT9), .B(KEYINPUT85), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U436 ( .A(G29GAT), .B(G134GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n377), .B(KEYINPUT86), .ZN(n410) );
  XNOR2_X1 U438 ( .A(n410), .B(n378), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n381), .B(G162GAT), .ZN(n383) );
  XOR2_X1 U441 ( .A(n387), .B(n386), .Z(n564) );
  INV_X1 U442 ( .A(n564), .ZN(n465) );
  NOR2_X1 U443 ( .A1(n576), .A2(n465), .ZN(n388) );
  NAND2_X1 U444 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n390), .B(KEYINPUT47), .ZN(n398) );
  INV_X1 U446 ( .A(n557), .ZN(n569) );
  XOR2_X1 U447 ( .A(KEYINPUT36), .B(KEYINPUT109), .Z(n391) );
  XNOR2_X1 U448 ( .A(n391), .B(n564), .ZN(n583) );
  INV_X1 U449 ( .A(n576), .ZN(n559) );
  NOR2_X1 U450 ( .A1(n583), .A2(n559), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n392), .B(KEYINPUT45), .ZN(n395) );
  INV_X1 U452 ( .A(n393), .ZN(n394) );
  NAND2_X1 U453 ( .A1(n395), .A2(n394), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n569), .A2(n396), .ZN(n397) );
  NOR2_X1 U455 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT48), .ZN(n532) );
  NOR2_X1 U457 ( .A1(n523), .A2(n532), .ZN(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT54), .B(n400), .ZN(n421) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT2), .Z(n402) );
  XNOR2_X1 U460 ( .A(G162GAT), .B(KEYINPUT96), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U462 ( .A(n403), .B(KEYINPUT3), .Z(n405) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(G155GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n429) );
  XOR2_X1 U465 ( .A(KEYINPUT4), .B(KEYINPUT100), .Z(n407) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U468 ( .A(n408), .B(KEYINPUT1), .Z(n412) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U471 ( .A(KEYINPUT6), .B(KEYINPUT101), .Z(n414) );
  XNOR2_X1 U472 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U474 ( .A(n416), .B(n415), .Z(n419) );
  XOR2_X1 U475 ( .A(G113GAT), .B(KEYINPUT0), .Z(n441) );
  XNOR2_X1 U476 ( .A(n441), .B(n417), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n429), .B(n420), .Z(n479) );
  XNOR2_X1 U479 ( .A(KEYINPUT102), .B(n479), .ZN(n521) );
  NAND2_X1 U480 ( .A1(n421), .A2(n521), .ZN(n423) );
  INV_X1 U481 ( .A(n568), .ZN(n439) );
  XOR2_X1 U482 ( .A(G148GAT), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U485 ( .A(n428), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U486 ( .A(G22GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(KEYINPUT98), .Z(n433) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U491 ( .A(n435), .B(n434), .Z(n438) );
  XNOR2_X1 U492 ( .A(n436), .B(KEYINPUT99), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n473) );
  XNOR2_X1 U494 ( .A(n440), .B(KEYINPUT55), .ZN(n460) );
  XOR2_X1 U495 ( .A(n441), .B(KEYINPUT65), .Z(n443) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n444), .B(G99GAT), .Z(n449) );
  XOR2_X1 U499 ( .A(KEYINPUT94), .B(KEYINPUT91), .Z(n446) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(KEYINPUT93), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U504 ( .A(G127GAT), .B(G190GAT), .Z(n451) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(G134GAT), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U507 ( .A(n453), .B(n452), .Z(n459) );
  XOR2_X1 U508 ( .A(G183GAT), .B(G176GAT), .Z(n455) );
  XNOR2_X1 U509 ( .A(KEYINPUT20), .B(G71GAT), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n533) );
  NOR2_X1 U513 ( .A1(n460), .A2(n533), .ZN(n461) );
  XNOR2_X1 U514 ( .A(KEYINPUT121), .B(n461), .ZN(n563) );
  NOR2_X1 U515 ( .A1(n548), .A2(n563), .ZN(n464) );
  XNOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n557), .A2(n393), .ZN(n498) );
  NOR2_X1 U518 ( .A1(n465), .A2(n559), .ZN(n466) );
  XNOR2_X1 U519 ( .A(KEYINPUT16), .B(n466), .ZN(n483) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(KEYINPUT103), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(n523), .ZN(n475) );
  INV_X1 U522 ( .A(n475), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n468), .A2(n521), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT104), .B(n469), .Z(n545) );
  XNOR2_X1 U525 ( .A(n473), .B(KEYINPUT28), .ZN(n491) );
  NOR2_X1 U526 ( .A1(n545), .A2(n491), .ZN(n535) );
  NAND2_X1 U527 ( .A1(n535), .A2(n533), .ZN(n481) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(KEYINPUT105), .Z(n472) );
  NOR2_X1 U529 ( .A1(n533), .A2(n523), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n473), .A2(n470), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n477) );
  NAND2_X1 U532 ( .A1(n473), .A2(n533), .ZN(n474) );
  XOR2_X1 U533 ( .A(n474), .B(KEYINPUT26), .Z(n567) );
  NAND2_X1 U534 ( .A1(n475), .A2(n567), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U538 ( .A(KEYINPUT106), .B(n482), .ZN(n495) );
  AND2_X1 U539 ( .A1(n483), .A2(n495), .ZN(n509) );
  NAND2_X1 U540 ( .A1(n498), .A2(n509), .ZN(n492) );
  NOR2_X1 U541 ( .A1(n521), .A2(n492), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(n484), .Z(n485) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n523), .A2(n492), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n533), .A2(n492), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT108), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n491), .ZN(n529) );
  NOR2_X1 U552 ( .A1(n529), .A2(n492), .ZN(n493) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n493), .Z(G1327GAT) );
  NOR2_X1 U554 ( .A1(n583), .A2(n576), .ZN(n494) );
  NAND2_X1 U555 ( .A1(n495), .A2(n494), .ZN(n497) );
  NAND2_X1 U556 ( .A1(n519), .A2(n498), .ZN(n499) );
  NOR2_X1 U557 ( .A1(n507), .A2(n521), .ZN(n501) );
  XNOR2_X1 U558 ( .A(KEYINPUT111), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U560 ( .A(G29GAT), .B(n502), .Z(G1328GAT) );
  NOR2_X1 U561 ( .A1(n507), .A2(n523), .ZN(n503) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  XNOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT112), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n533), .A2(n507), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U566 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U567 ( .A1(n529), .A2(n507), .ZN(n508) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NOR2_X1 U569 ( .A1(n548), .A2(n569), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n520), .A2(n509), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n521), .A2(n515), .ZN(n511) );
  XNOR2_X1 U572 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n523), .A2(n515), .ZN(n513) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n533), .A2(n515), .ZN(n514) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n529), .A2(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n521), .A2(n528), .ZN(n522) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n528), .ZN(n525) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n533), .A2(n528), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT116), .B(n526), .Z(n527) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n542) );
  NOR2_X1 U597 ( .A1(n557), .A2(n542), .ZN(n536) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n548), .A2(n542), .ZN(n538) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n559), .A2(n542), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  NOR2_X1 U606 ( .A1(n564), .A2(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n545), .A2(n532), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n546), .A2(n567), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n557), .A2(n553), .ZN(n547) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n553), .ZN(n550) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n559), .A2(n553), .ZN(n552) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n564), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n558) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n563), .ZN(n560) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n562) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n566) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(n566), .B(n565), .Z(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n582) );
  INV_X1 U634 ( .A(n582), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U639 ( .A1(n577), .A2(n393), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

