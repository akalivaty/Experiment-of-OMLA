

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754;

  BUF_X1 U371 ( .A(n623), .Z(n350) );
  XNOR2_X1 U372 ( .A(n516), .B(KEYINPUT101), .ZN(n749) );
  NAND2_X1 U373 ( .A1(n370), .A2(n368), .ZN(n516) );
  AND2_X1 U374 ( .A1(n355), .A2(n351), .ZN(n542) );
  BUF_X1 U375 ( .A(n518), .Z(n669) );
  INV_X1 U376 ( .A(n563), .ZN(n512) );
  NAND2_X1 U377 ( .A1(n380), .A2(n376), .ZN(n540) );
  XOR2_X1 U378 ( .A(G140), .B(KEYINPUT70), .Z(n466) );
  XNOR2_X1 U379 ( .A(G107), .B(G104), .ZN(n464) );
  INV_X1 U380 ( .A(G128), .ZN(n430) );
  INV_X1 U381 ( .A(KEYINPUT64), .ZN(n425) );
  NOR2_X2 U382 ( .A1(n584), .A2(n521), .ZN(n351) );
  INV_X1 U383 ( .A(n539), .ZN(n535) );
  XNOR2_X2 U384 ( .A(n597), .B(n596), .ZN(n730) );
  XNOR2_X2 U385 ( .A(n736), .B(n471), .ZN(n707) );
  XNOR2_X1 U386 ( .A(G101), .B(G110), .ZN(n465) );
  NAND2_X1 U387 ( .A1(n527), .A2(n669), .ZN(n528) );
  XNOR2_X1 U388 ( .A(n475), .B(n476), .ZN(n477) );
  XNOR2_X2 U389 ( .A(n536), .B(n504), .ZN(n636) );
  NAND2_X2 U390 ( .A1(n580), .A2(n579), .ZN(n364) );
  NAND2_X2 U391 ( .A1(n608), .A2(n660), .ZN(n610) );
  AND2_X1 U392 ( .A1(n374), .A2(n371), .ZN(n370) );
  NOR2_X1 U393 ( .A1(n685), .A2(n684), .ZN(n398) );
  NOR2_X1 U394 ( .A1(n563), .A2(n666), .ZN(n663) );
  AND2_X1 U395 ( .A1(n382), .A2(n381), .ZN(n380) );
  OR2_X1 U396 ( .A1(n611), .A2(n377), .ZN(n376) );
  XNOR2_X1 U397 ( .A(n409), .B(n408), .ZN(n611) );
  NAND2_X1 U398 ( .A1(n707), .A2(n378), .ZN(n474) );
  NOR2_X1 U399 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U400 ( .A(n396), .B(n395), .ZN(n754) );
  NOR2_X1 U401 ( .A1(n586), .A2(n669), .ZN(n638) );
  NAND2_X1 U402 ( .A1(n369), .A2(KEYINPUT36), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n398), .B(n530), .ZN(n699) );
  NAND2_X1 U404 ( .A1(n457), .A2(n680), .ZN(n514) );
  NAND2_X1 U405 ( .A1(n385), .A2(n383), .ZN(n539) );
  XOR2_X1 U406 ( .A(KEYINPUT121), .B(n611), .Z(n612) );
  NAND2_X1 U407 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X1 U408 ( .A(G137), .B(KEYINPUT68), .ZN(n480) );
  XNOR2_X1 U409 ( .A(n499), .B(n498), .ZN(n630) );
  XNOR2_X1 U410 ( .A(n364), .B(n581), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n364), .B(n581), .ZN(n747) );
  XNOR2_X2 U412 ( .A(n459), .B(KEYINPUT0), .ZN(n587) );
  XOR2_X1 U413 ( .A(KEYINPUT59), .B(n350), .Z(n624) );
  XNOR2_X1 U414 ( .A(n423), .B(n422), .ZN(n623) );
  XNOR2_X2 U415 ( .A(n525), .B(KEYINPUT40), .ZN(n752) );
  AND2_X1 U416 ( .A1(n534), .A2(n533), .ZN(n649) );
  XNOR2_X1 U417 ( .A(n393), .B(n356), .ZN(n725) );
  XNOR2_X2 U418 ( .A(n501), .B(n500), .ZN(n518) );
  XNOR2_X2 U419 ( .A(n417), .B(KEYINPUT10), .ZN(n481) );
  XNOR2_X2 U420 ( .A(G125), .B(G140), .ZN(n417) );
  XNOR2_X2 U421 ( .A(KEYINPUT4), .B(G146), .ZN(n461) );
  OR2_X1 U422 ( .A1(n543), .A2(n648), .ZN(n544) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n490) );
  INV_X1 U424 ( .A(n599), .ZN(n406) );
  INV_X1 U425 ( .A(KEYINPUT67), .ZN(n405) );
  NAND2_X1 U426 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U427 ( .A(n560), .B(n559), .ZN(n603) );
  NAND2_X1 U428 ( .A1(n558), .A2(n659), .ZN(n560) );
  NAND2_X1 U429 ( .A1(n611), .A2(G478), .ZN(n382) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n456) );
  AND2_X1 U431 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U432 ( .A1(n424), .A2(n378), .ZN(n384) );
  BUF_X1 U433 ( .A(n573), .Z(n662) );
  XNOR2_X1 U434 ( .A(n445), .B(KEYINPUT16), .ZN(n394) );
  XNOR2_X1 U435 ( .A(G146), .B(G128), .ZN(n476) );
  INV_X1 U436 ( .A(KEYINPUT24), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n427), .B(n426), .ZN(n478) );
  INV_X1 U438 ( .A(KEYINPUT8), .ZN(n426) );
  XNOR2_X1 U439 ( .A(n428), .B(n412), .ZN(n411) );
  XOR2_X1 U440 ( .A(G143), .B(G131), .Z(n420) );
  XNOR2_X1 U441 ( .A(G113), .B(G146), .ZN(n419) );
  XNOR2_X1 U442 ( .A(n481), .B(KEYINPUT12), .ZN(n360) );
  XOR2_X1 U443 ( .A(KEYINPUT91), .B(KEYINPUT11), .Z(n416) );
  XNOR2_X1 U444 ( .A(n725), .B(n389), .ZN(n617) );
  XNOR2_X1 U445 ( .A(n453), .B(n390), .ZN(n389) );
  NAND2_X1 U446 ( .A1(n363), .A2(n362), .ZN(n460) );
  NOR2_X1 U447 ( .A1(n684), .A2(n666), .ZN(n362) );
  NOR2_X1 U448 ( .A1(n397), .A2(n529), .ZN(n534) );
  XNOR2_X1 U449 ( .A(n528), .B(KEYINPUT28), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n488), .B(n487), .ZN(n563) );
  NAND2_X1 U451 ( .A1(n388), .A2(G902), .ZN(n386) );
  NAND2_X1 U452 ( .A1(n406), .A2(n405), .ZN(n404) );
  NOR2_X1 U453 ( .A1(n403), .A2(n402), .ZN(n401) );
  AND2_X1 U454 ( .A1(n599), .A2(KEYINPUT2), .ZN(n403) );
  NOR2_X1 U455 ( .A1(n602), .A2(n405), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n461), .B(n392), .ZN(n391) );
  INV_X1 U457 ( .A(KEYINPUT70), .ZN(n392) );
  XNOR2_X1 U458 ( .A(G125), .B(KEYINPUT82), .ZN(n449) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n450) );
  INV_X1 U460 ( .A(G478), .ZN(n379) );
  NAND2_X1 U461 ( .A1(G902), .A2(G478), .ZN(n381) );
  XNOR2_X1 U462 ( .A(G902), .B(KEYINPUT15), .ZN(n601) );
  XOR2_X1 U463 ( .A(G119), .B(KEYINPUT5), .Z(n492) );
  XNOR2_X1 U464 ( .A(KEYINPUT89), .B(G137), .ZN(n493) );
  XNOR2_X1 U465 ( .A(n695), .B(n694), .ZN(n696) );
  AND2_X1 U466 ( .A1(n372), .A2(n662), .ZN(n371) );
  NAND2_X1 U467 ( .A1(n373), .A2(KEYINPUT36), .ZN(n372) );
  INV_X1 U468 ( .A(n515), .ZN(n373) );
  XNOR2_X1 U469 ( .A(n514), .B(KEYINPUT19), .ZN(n533) );
  INV_X1 U470 ( .A(KEYINPUT97), .ZN(n504) );
  XNOR2_X1 U471 ( .A(n394), .B(n496), .ZN(n393) );
  XNOR2_X1 U472 ( .A(n479), .B(n365), .ZN(n483) );
  XNOR2_X1 U473 ( .A(n477), .B(n366), .ZN(n365) );
  NAND2_X1 U474 ( .A1(n478), .A2(G217), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n360), .B(n418), .ZN(n423) );
  INV_X1 U476 ( .A(KEYINPUT42), .ZN(n395) );
  NAND2_X1 U477 ( .A1(n699), .A2(n534), .ZN(n396) );
  INV_X1 U478 ( .A(KEYINPUT32), .ZN(n571) );
  NOR2_X1 U479 ( .A1(n503), .A2(n502), .ZN(n592) );
  AND2_X1 U480 ( .A1(n603), .A2(n358), .ZN(n353) );
  AND2_X1 U481 ( .A1(n701), .A2(n414), .ZN(n354) );
  XOR2_X1 U482 ( .A(KEYINPUT30), .B(n519), .Z(n355) );
  XOR2_X1 U483 ( .A(n447), .B(n475), .Z(n356) );
  AND2_X1 U484 ( .A1(n607), .A2(n658), .ZN(n357) );
  AND2_X1 U485 ( .A1(n658), .A2(n404), .ZN(n358) );
  AND2_X1 U486 ( .A1(n515), .A2(n400), .ZN(n359) );
  INV_X1 U487 ( .A(G902), .ZN(n378) );
  INV_X1 U488 ( .A(KEYINPUT36), .ZN(n400) );
  NAND2_X1 U489 ( .A1(n595), .A2(n361), .ZN(n597) );
  XNOR2_X1 U490 ( .A(n583), .B(KEYINPUT44), .ZN(n361) );
  INV_X1 U491 ( .A(n730), .ZN(n598) );
  NAND2_X1 U492 ( .A1(n747), .A2(n751), .ZN(n582) );
  NOR2_X1 U493 ( .A1(n689), .A2(n587), .ZN(n577) );
  XNOR2_X1 U494 ( .A(n526), .B(KEYINPUT1), .ZN(n573) );
  NAND2_X1 U495 ( .A1(n533), .A2(n458), .ZN(n459) );
  NOR2_X2 U496 ( .A1(n582), .A2(n643), .ZN(n583) );
  INV_X1 U497 ( .A(n587), .ZN(n363) );
  NOR2_X1 U498 ( .A1(n717), .A2(n722), .ZN(G54) );
  XNOR2_X1 U499 ( .A(n367), .B(n391), .ZN(n390) );
  XNOR2_X2 U500 ( .A(n367), .B(G134), .ZN(n463) );
  XNOR2_X2 U501 ( .A(n431), .B(n430), .ZN(n367) );
  INV_X1 U502 ( .A(n375), .ZN(n369) );
  NAND2_X1 U503 ( .A1(n375), .A2(n359), .ZN(n374) );
  XNOR2_X1 U504 ( .A(n550), .B(KEYINPUT100), .ZN(n375) );
  NOR2_X4 U505 ( .A1(n535), .A2(n540), .ZN(n536) );
  OR2_X1 U506 ( .A1(n623), .A2(n384), .ZN(n383) );
  NAND2_X1 U507 ( .A1(n623), .A2(n388), .ZN(n387) );
  INV_X1 U508 ( .A(n424), .ZN(n388) );
  XNOR2_X2 U509 ( .A(n448), .B(G101), .ZN(n496) );
  XNOR2_X2 U510 ( .A(KEYINPUT22), .B(n460), .ZN(n570) );
  NOR2_X2 U511 ( .A1(n512), .A2(n511), .ZN(n527) );
  NAND2_X1 U512 ( .A1(n399), .A2(n401), .ZN(n608) );
  NAND2_X1 U513 ( .A1(n598), .A2(n353), .ZN(n399) );
  NAND2_X1 U514 ( .A1(n598), .A2(n357), .ZN(n407) );
  NAND2_X1 U515 ( .A1(n407), .A2(n600), .ZN(n661) );
  XNOR2_X1 U516 ( .A(n463), .B(n410), .ZN(n409) );
  XNOR2_X1 U517 ( .A(n413), .B(n411), .ZN(n410) );
  INV_X1 U518 ( .A(KEYINPUT93), .ZN(n412) );
  XNOR2_X1 U519 ( .A(n429), .B(n446), .ZN(n413) );
  NOR2_X2 U520 ( .A1(n570), .A2(n662), .ZN(n562) );
  NOR2_X2 U521 ( .A1(n570), .A2(n569), .ZN(n572) );
  BUF_X1 U522 ( .A(n636), .Z(n651) );
  OR2_X1 U523 ( .A1(n700), .A2(n690), .ZN(n414) );
  XNOR2_X1 U524 ( .A(n668), .B(KEYINPUT49), .ZN(n670) );
  XNOR2_X1 U525 ( .A(n675), .B(KEYINPUT110), .ZN(n676) );
  XNOR2_X1 U526 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U527 ( .A(KEYINPUT114), .B(KEYINPUT52), .ZN(n694) );
  INV_X1 U528 ( .A(n520), .ZN(n521) );
  OR2_X1 U529 ( .A1(n742), .A2(G952), .ZN(n633) );
  INV_X1 U530 ( .A(n752), .ZN(n753) );
  NAND2_X1 U531 ( .A1(G214), .A2(n490), .ZN(n415) );
  XNOR2_X1 U532 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X2 U533 ( .A(G122), .B(G104), .ZN(n444) );
  XNOR2_X1 U534 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U535 ( .A(n444), .B(n421), .ZN(n422) );
  XNOR2_X1 U536 ( .A(KEYINPUT13), .B(G475), .ZN(n424) );
  XNOR2_X2 U537 ( .A(n425), .B(G953), .ZN(n742) );
  NAND2_X1 U538 ( .A1(n742), .A2(G234), .ZN(n427) );
  XNOR2_X1 U539 ( .A(G116), .B(G107), .ZN(n446) );
  XOR2_X1 U540 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n429) );
  XNOR2_X1 U541 ( .A(G122), .B(KEYINPUT92), .ZN(n428) );
  XNOR2_X2 U542 ( .A(KEYINPUT76), .B(G143), .ZN(n431) );
  INV_X1 U543 ( .A(n540), .ZN(n432) );
  NAND2_X1 U544 ( .A1(n535), .A2(n432), .ZN(n684) );
  XOR2_X1 U545 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n436) );
  XOR2_X1 U546 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n434) );
  NAND2_X1 U547 ( .A1(G234), .A2(n601), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n434), .B(n433), .ZN(n484) );
  NAND2_X1 U549 ( .A1(G221), .A2(n484), .ZN(n435) );
  XNOR2_X1 U550 ( .A(n436), .B(n435), .ZN(n666) );
  XNOR2_X1 U551 ( .A(n437), .B(KEYINPUT14), .ZN(n438) );
  XNOR2_X1 U552 ( .A(KEYINPUT72), .B(n438), .ZN(n441) );
  NAND2_X1 U553 ( .A1(G902), .A2(n441), .ZN(n505) );
  INV_X1 U554 ( .A(n505), .ZN(n439) );
  INV_X1 U555 ( .A(G953), .ZN(n739) );
  NOR2_X1 U556 ( .A1(G898), .A2(n739), .ZN(n726) );
  NAND2_X1 U557 ( .A1(n439), .A2(n726), .ZN(n440) );
  XNOR2_X1 U558 ( .A(n440), .B(KEYINPUT84), .ZN(n443) );
  NAND2_X1 U559 ( .A1(G952), .A2(n441), .ZN(n697) );
  NOR2_X1 U560 ( .A1(G953), .A2(n697), .ZN(n442) );
  XNOR2_X1 U561 ( .A(KEYINPUT83), .B(n442), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n443), .A2(n509), .ZN(n458) );
  INV_X1 U563 ( .A(n444), .ZN(n445) );
  INV_X1 U564 ( .A(n446), .ZN(n447) );
  XOR2_X2 U565 ( .A(G119), .B(G110), .Z(n475) );
  XNOR2_X2 U566 ( .A(KEYINPUT3), .B(G113), .ZN(n448) );
  XNOR2_X1 U567 ( .A(n450), .B(n449), .ZN(n452) );
  NAND2_X1 U568 ( .A1(n742), .A2(G224), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U570 ( .A1(n617), .A2(n601), .ZN(n455) );
  NAND2_X1 U571 ( .A1(G210), .A2(n456), .ZN(n454) );
  XNOR2_X2 U572 ( .A(n455), .B(n454), .ZN(n556) );
  INV_X1 U573 ( .A(n556), .ZN(n457) );
  NAND2_X1 U574 ( .A1(n456), .A2(G214), .ZN(n680) );
  XNOR2_X1 U575 ( .A(n461), .B(G131), .ZN(n462) );
  XNOR2_X2 U576 ( .A(n463), .B(n462), .ZN(n736) );
  XNOR2_X1 U577 ( .A(n464), .B(n480), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n468), .B(n467), .ZN(n470) );
  NAND2_X1 U580 ( .A1(G227), .A2(n742), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n470), .B(n469), .ZN(n471) );
  INV_X1 U582 ( .A(KEYINPUT69), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n472), .B(G469), .ZN(n473) );
  XNOR2_X2 U584 ( .A(n474), .B(n473), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n478), .A2(G221), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n735) );
  XNOR2_X1 U587 ( .A(n735), .B(KEYINPUT23), .ZN(n482) );
  XNOR2_X1 U588 ( .A(n483), .B(n482), .ZN(n719) );
  NOR2_X1 U589 ( .A1(n719), .A2(G902), .ZN(n488) );
  XOR2_X1 U590 ( .A(KEYINPUT86), .B(KEYINPUT25), .Z(n486) );
  NAND2_X1 U591 ( .A1(n484), .A2(G217), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U593 ( .A(n512), .B(KEYINPUT94), .Z(n667) );
  INV_X1 U594 ( .A(n667), .ZN(n489) );
  NAND2_X1 U595 ( .A1(n562), .A2(n489), .ZN(n503) );
  INV_X1 U596 ( .A(n736), .ZN(n499) );
  NAND2_X1 U597 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n492), .B(n491), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n493), .B(G116), .ZN(n494) );
  XNOR2_X1 U600 ( .A(n495), .B(n494), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X2 U602 ( .A1(n630), .A2(G902), .ZN(n501) );
  XOR2_X1 U603 ( .A(G472), .B(KEYINPUT90), .Z(n500) );
  XNOR2_X1 U604 ( .A(n518), .B(KEYINPUT6), .ZN(n574) );
  INV_X1 U605 ( .A(n574), .ZN(n502) );
  XOR2_X1 U606 ( .A(G101), .B(n592), .Z(G3) );
  INV_X1 U607 ( .A(n666), .ZN(n510) );
  NOR2_X1 U608 ( .A1(G900), .A2(n505), .ZN(n507) );
  INV_X1 U609 ( .A(n742), .ZN(n506) );
  NAND2_X1 U610 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U611 ( .A1(n509), .A2(n508), .ZN(n520) );
  NAND2_X1 U612 ( .A1(n510), .A2(n520), .ZN(n511) );
  NAND2_X1 U613 ( .A1(n636), .A2(n527), .ZN(n513) );
  NOR2_X2 U614 ( .A1(n513), .A2(n574), .ZN(n550) );
  INV_X1 U615 ( .A(n514), .ZN(n515) );
  INV_X1 U616 ( .A(KEYINPUT80), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n749), .B(n517), .ZN(n547) );
  NAND2_X1 U618 ( .A1(n518), .A2(n680), .ZN(n519) );
  NAND2_X1 U619 ( .A1(n526), .A2(n663), .ZN(n584) );
  XNOR2_X1 U620 ( .A(KEYINPUT38), .B(n556), .ZN(n681) );
  NAND2_X1 U621 ( .A1(n542), .A2(n681), .ZN(n524) );
  XOR2_X1 U622 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n523) );
  XNOR2_X1 U623 ( .A(n524), .B(n523), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n561), .A2(n536), .ZN(n525) );
  INV_X1 U625 ( .A(n526), .ZN(n529) );
  NAND2_X1 U626 ( .A1(n681), .A2(n680), .ZN(n685) );
  XNOR2_X1 U627 ( .A(KEYINPUT99), .B(KEYINPUT41), .ZN(n530) );
  INV_X1 U628 ( .A(n754), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n752), .A2(n531), .ZN(n532) );
  XNOR2_X1 U630 ( .A(n532), .B(KEYINPUT46), .ZN(n545) );
  AND2_X1 U631 ( .A1(n540), .A2(n535), .ZN(n654) );
  NOR2_X1 U632 ( .A1(n536), .A2(n654), .ZN(n686) );
  INV_X1 U633 ( .A(n686), .ZN(n537) );
  NAND2_X1 U634 ( .A1(n649), .A2(n537), .ZN(n538) );
  XNOR2_X1 U635 ( .A(n538), .B(KEYINPUT47), .ZN(n543) );
  NAND2_X1 U636 ( .A1(n540), .A2(n539), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n578), .A2(n556), .ZN(n541) );
  AND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n648) );
  NAND2_X1 U639 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U640 ( .A(KEYINPUT79), .B(KEYINPUT48), .ZN(n548) );
  XNOR2_X1 U641 ( .A(n549), .B(n548), .ZN(n558) );
  BUF_X1 U642 ( .A(n550), .Z(n553) );
  INV_X1 U643 ( .A(n680), .ZN(n551) );
  NOR2_X1 U644 ( .A1(n662), .A2(n551), .ZN(n552) );
  NAND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U646 ( .A(KEYINPUT43), .B(KEYINPUT98), .ZN(n554) );
  XNOR2_X1 U647 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n659) );
  INV_X1 U649 ( .A(KEYINPUT78), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n561), .A2(n654), .ZN(n658) );
  INV_X1 U651 ( .A(n562), .ZN(n565) );
  INV_X1 U652 ( .A(n669), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n563), .A2(n588), .ZN(n564) );
  NOR2_X1 U654 ( .A1(n565), .A2(n564), .ZN(n643) );
  NAND2_X1 U655 ( .A1(n667), .A2(n574), .ZN(n567) );
  INV_X1 U656 ( .A(n662), .ZN(n566) );
  NOR2_X1 U657 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U658 ( .A(n568), .B(KEYINPUT75), .ZN(n569) );
  XNOR2_X2 U659 ( .A(n572), .B(n571), .ZN(n751) );
  XNOR2_X1 U660 ( .A(KEYINPUT73), .B(KEYINPUT35), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n573), .A2(n663), .ZN(n589) );
  XNOR2_X1 U662 ( .A(KEYINPUT96), .B(n589), .ZN(n575) );
  NOR2_X1 U663 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U664 ( .A(n576), .B(KEYINPUT33), .ZN(n689) );
  XNOR2_X1 U665 ( .A(n577), .B(KEYINPUT34), .ZN(n580) );
  XOR2_X1 U666 ( .A(n578), .B(KEYINPUT74), .Z(n579) );
  NOR2_X1 U667 ( .A1(n587), .A2(n584), .ZN(n585) );
  XOR2_X1 U668 ( .A(KEYINPUT88), .B(n585), .Z(n586) );
  NOR2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n673) );
  NAND2_X1 U670 ( .A1(n363), .A2(n673), .ZN(n590) );
  XNOR2_X1 U671 ( .A(n590), .B(KEYINPUT31), .ZN(n655) );
  NOR2_X1 U672 ( .A1(n638), .A2(n655), .ZN(n591) );
  NOR2_X1 U673 ( .A1(n591), .A2(n686), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U675 ( .A(KEYINPUT95), .B(n594), .Z(n595) );
  XNOR2_X1 U676 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n596) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(KEYINPUT67), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n602) );
  BUF_X1 U680 ( .A(n603), .Z(n607) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(n658), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT77), .B(n604), .Z(n605) );
  NOR2_X1 U683 ( .A1(n730), .A2(n605), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n660) );
  INV_X1 U685 ( .A(KEYINPUT66), .ZN(n609) );
  XNOR2_X2 U686 ( .A(n610), .B(n609), .ZN(n718) );
  NAND2_X1 U687 ( .A1(n718), .A2(G478), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(n614) );
  INV_X1 U689 ( .A(n633), .ZN(n722) );
  NOR2_X2 U690 ( .A1(n614), .A2(n722), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U692 ( .A1(n718), .A2(G210), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U696 ( .A1(n620), .A2(n722), .ZN(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT118), .B(KEYINPUT56), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(G51) );
  NAND2_X1 U699 ( .A1(n718), .A2(G475), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U701 ( .A1(n626), .A2(n722), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U703 ( .A1(n718), .A2(G472), .ZN(n632) );
  XNOR2_X1 U704 ( .A(KEYINPUT81), .B(KEYINPUT102), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT62), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n632), .B(n631), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n635), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n638), .A2(n651), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(G104), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U713 ( .A1(n638), .A2(n654), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n642) );
  XOR2_X1 U715 ( .A(G107), .B(KEYINPUT103), .Z(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(G9) );
  XOR2_X1 U717 ( .A(G110), .B(n643), .Z(G12) );
  XOR2_X1 U718 ( .A(KEYINPUT105), .B(KEYINPUT29), .Z(n645) );
  NAND2_X1 U719 ( .A1(n649), .A2(n654), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(n647) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT104), .Z(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(G30) );
  XOR2_X1 U723 ( .A(G143), .B(n648), .Z(G45) );
  NAND2_X1 U724 ( .A1(n651), .A2(n649), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(G146), .ZN(G48) );
  NAND2_X1 U726 ( .A1(n655), .A2(n651), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n652), .B(KEYINPUT106), .ZN(n653) );
  XNOR2_X1 U728 ( .A(G113), .B(n653), .ZN(G15) );
  XOR2_X1 U729 ( .A(G116), .B(KEYINPUT107), .Z(n657) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n657), .B(n656), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G134), .B(n658), .ZN(G36) );
  XNOR2_X1 U733 ( .A(G140), .B(n659), .ZN(G42) );
  AND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n703) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT50), .B(KEYINPUT109), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  AND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n677) );
  XOR2_X1 U742 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n675) );
  NAND2_X1 U743 ( .A1(n699), .A2(n678), .ZN(n679) );
  XOR2_X1 U744 ( .A(KEYINPUT112), .B(n679), .Z(n693) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT113), .B(n682), .Z(n683) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n691) );
  BUF_X1 U750 ( .A(n689), .Z(n690) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT115), .ZN(n701) );
  INV_X1 U755 ( .A(n699), .ZN(n700) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(n354), .Z(n702) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n704), .B(KEYINPUT117), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U760 ( .A(KEYINPUT53), .B(n706), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n718), .A2(G469), .ZN(n710) );
  INV_X1 U762 ( .A(n710), .ZN(n709) );
  INV_X1 U763 ( .A(n707), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n710), .A2(n707), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n716) );
  XOR2_X1 U767 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n714) );
  XNOR2_X1 U768 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U771 ( .A1(n718), .A2(G217), .ZN(n721) );
  XOR2_X1 U772 ( .A(n719), .B(KEYINPUT123), .Z(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n723) );
  NOR2_X2 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n724), .B(KEYINPUT124), .ZN(G66) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n734) );
  XOR2_X1 U777 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n728) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n729), .A2(G898), .ZN(n732) );
  OR2_X1 U781 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(G69) );
  XOR2_X1 U784 ( .A(n736), .B(n735), .Z(n741) );
  XOR2_X1 U785 ( .A(G227), .B(n741), .Z(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G900), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(KEYINPUT126), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G953), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n357), .B(n741), .ZN(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n745), .A2(n744), .ZN(G72) );
  XOR2_X1 U792 ( .A(G122), .B(KEYINPUT127), .Z(n746) );
  XNOR2_X1 U793 ( .A(n352), .B(n746), .ZN(G24) );
  XNOR2_X1 U794 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n748) );
  XNOR2_X1 U795 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U796 ( .A(G125), .B(n750), .ZN(G27) );
  XNOR2_X1 U797 ( .A(G119), .B(n751), .ZN(G21) );
  XOR2_X1 U798 ( .A(G131), .B(n753), .Z(G33) );
  XOR2_X1 U799 ( .A(G137), .B(n754), .Z(G39) );
endmodule

