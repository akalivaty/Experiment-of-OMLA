

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n687), .A2(n515), .ZN(n688) );
  NAND2_X1 U551 ( .A1(n683), .A2(n741), .ZN(n722) );
  NOR2_X1 U552 ( .A1(G164), .A2(G1384), .ZN(n741) );
  XNOR2_X1 U553 ( .A(n518), .B(KEYINPUT65), .ZN(n870) );
  AND2_X1 U554 ( .A1(n722), .A2(G1341), .ZN(n515) );
  XOR2_X1 U555 ( .A(KEYINPUT99), .B(n713), .Z(n516) );
  XOR2_X1 U556 ( .A(n721), .B(KEYINPUT31), .Z(n517) );
  INV_X1 U557 ( .A(KEYINPUT27), .ZN(n695) );
  INV_X1 U558 ( .A(n722), .ZN(n708) );
  NOR2_X1 U559 ( .A1(n694), .A2(n693), .ZN(n701) );
  NOR2_X1 U560 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U561 ( .A1(n516), .A2(n517), .ZN(n733) );
  AND2_X1 U562 ( .A1(n680), .A2(G40), .ZN(n681) );
  XNOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n730) );
  NAND2_X1 U564 ( .A1(n682), .A2(n681), .ZN(n740) );
  XOR2_X1 U565 ( .A(KEYINPUT64), .B(G2104), .Z(n522) );
  NOR2_X2 U566 ( .A1(n522), .A2(G2105), .ZN(n876) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n519), .Z(n875) );
  NOR2_X1 U568 ( .A1(G651), .A2(n625), .ZN(n651) );
  NAND2_X1 U569 ( .A1(G2105), .A2(n522), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n870), .A2(G126), .ZN(n521) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  NAND2_X1 U572 ( .A1(n875), .A2(G138), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n526) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U575 ( .A1(G114), .A2(n871), .ZN(n524) );
  NAND2_X1 U576 ( .A1(G102), .A2(n876), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(G164) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U580 ( .A1(n642), .A2(G89), .ZN(n527) );
  XNOR2_X1 U581 ( .A(n527), .B(KEYINPUT4), .ZN(n529) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n625) );
  INV_X1 U583 ( .A(G651), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n625), .A2(n531), .ZN(n646) );
  NAND2_X1 U585 ( .A1(G76), .A2(n646), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n530), .B(KEYINPUT5), .ZN(n538) );
  XNOR2_X1 U588 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G51), .A2(n651), .ZN(n534) );
  NOR2_X1 U590 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n532), .Z(n640) );
  NAND2_X1 U592 ( .A1(G63), .A2(n640), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U594 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(KEYINPUT7), .B(n539), .ZN(G168) );
  XOR2_X1 U597 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U598 ( .A1(G53), .A2(n651), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G65), .A2(n640), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G78), .A2(n646), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G91), .A2(n642), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U604 ( .A(KEYINPUT70), .B(n544), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U606 ( .A(n547), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U607 ( .A1(G125), .A2(n870), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G137), .A2(n875), .ZN(n549) );
  NAND2_X1 U609 ( .A1(G113), .A2(n871), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT67), .ZN(n551) );
  AND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n682) );
  NAND2_X1 U613 ( .A1(G101), .A2(n876), .ZN(n553) );
  XNOR2_X1 U614 ( .A(n553), .B(KEYINPUT23), .ZN(n554) );
  XOR2_X1 U615 ( .A(n554), .B(KEYINPUT66), .Z(n680) );
  AND2_X1 U616 ( .A1(n682), .A2(n680), .ZN(G160) );
  NAND2_X1 U617 ( .A1(G77), .A2(n646), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G90), .A2(n642), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G52), .A2(n651), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G64), .A2(n640), .ZN(n560) );
  XNOR2_X1 U624 ( .A(KEYINPUT69), .B(n560), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n562), .A2(n561), .ZN(G171) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  INV_X1 U628 ( .A(G132), .ZN(G219) );
  INV_X1 U629 ( .A(G82), .ZN(G220) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n565) );
  INV_X1 U633 ( .A(G223), .ZN(n826) );
  NAND2_X1 U634 ( .A1(G567), .A2(n826), .ZN(n564) );
  XNOR2_X1 U635 ( .A(n565), .B(n564), .ZN(G234) );
  NAND2_X1 U636 ( .A1(n651), .A2(G43), .ZN(n566) );
  XNOR2_X1 U637 ( .A(KEYINPUT76), .B(n566), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n640), .A2(G56), .ZN(n567) );
  XNOR2_X1 U639 ( .A(KEYINPUT14), .B(n567), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n569) );
  NAND2_X1 U641 ( .A1(G81), .A2(n642), .ZN(n568) );
  XNOR2_X1 U642 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U643 ( .A(KEYINPUT73), .B(n570), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n646), .A2(G68), .ZN(n571) );
  NAND2_X1 U645 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U646 ( .A(KEYINPUT13), .B(n573), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U648 ( .A(KEYINPUT75), .B(n576), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n955) );
  INV_X1 U650 ( .A(G860), .ZN(n592) );
  OR2_X1 U651 ( .A1(n955), .A2(n592), .ZN(G153) );
  XNOR2_X1 U652 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n579) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT78), .ZN(n588) );
  INV_X1 U655 ( .A(G868), .ZN(n664) );
  NAND2_X1 U656 ( .A1(G79), .A2(n646), .ZN(n581) );
  NAND2_X1 U657 ( .A1(G92), .A2(n642), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G54), .A2(n651), .ZN(n583) );
  NAND2_X1 U660 ( .A1(G66), .A2(n640), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT15), .ZN(n692) );
  NAND2_X1 U664 ( .A1(n664), .A2(n692), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(G284) );
  XNOR2_X1 U666 ( .A(KEYINPUT80), .B(n664), .ZN(n589) );
  NOR2_X1 U667 ( .A1(G286), .A2(n589), .ZN(n591) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n592), .A2(G559), .ZN(n593) );
  INV_X1 U671 ( .A(n692), .ZN(n958) );
  NAND2_X1 U672 ( .A1(n593), .A2(n958), .ZN(n594) );
  XNOR2_X1 U673 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G559), .A2(n664), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n958), .A2(n595), .ZN(n596) );
  XNOR2_X1 U676 ( .A(n596), .B(KEYINPUT81), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n955), .A2(G868), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G135), .A2(n875), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G111), .A2(n871), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n870), .A2(G123), .ZN(n601) );
  XNOR2_X1 U683 ( .A(n601), .B(KEYINPUT18), .ZN(n603) );
  NAND2_X1 U684 ( .A1(G99), .A2(n876), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n995) );
  XNOR2_X1 U687 ( .A(n995), .B(G2096), .ZN(n607) );
  INV_X1 U688 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G55), .A2(n651), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G67), .A2(n640), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G80), .A2(n646), .ZN(n611) );
  NAND2_X1 U694 ( .A1(G93), .A2(n642), .ZN(n610) );
  NAND2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n663) );
  XNOR2_X1 U697 ( .A(KEYINPUT82), .B(n955), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n958), .A2(G559), .ZN(n661) );
  XNOR2_X1 U699 ( .A(n614), .B(n661), .ZN(n615) );
  NOR2_X1 U700 ( .A1(G860), .A2(n615), .ZN(n616) );
  XOR2_X1 U701 ( .A(n663), .B(n616), .Z(G145) );
  NAND2_X1 U702 ( .A1(n640), .A2(G62), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G75), .A2(n646), .ZN(n618) );
  NAND2_X1 U704 ( .A1(G88), .A2(n642), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n651), .A2(G50), .ZN(n619) );
  XOR2_X1 U707 ( .A(KEYINPUT88), .B(n619), .Z(n620) );
  NOR2_X1 U708 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U710 ( .A(KEYINPUT89), .B(n624), .Z(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G87), .A2(n625), .ZN(n626) );
  XNOR2_X1 U713 ( .A(n626), .B(KEYINPUT84), .ZN(n629) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n627) );
  XOR2_X1 U715 ( .A(KEYINPUT83), .B(n627), .Z(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U717 ( .A1(n640), .A2(n630), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n651), .A2(G49), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G47), .A2(n651), .ZN(n634) );
  NAND2_X1 U721 ( .A1(G60), .A2(n640), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G72), .A2(n646), .ZN(n635) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(n635), .Z(n636) );
  NOR2_X1 U725 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n642), .A2(G85), .ZN(n638) );
  NAND2_X1 U727 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U728 ( .A1(n640), .A2(G61), .ZN(n641) );
  XOR2_X1 U729 ( .A(KEYINPUT85), .B(n641), .Z(n644) );
  NAND2_X1 U730 ( .A1(n642), .A2(G86), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U732 ( .A(KEYINPUT86), .B(n645), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U734 ( .A(n647), .B(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U735 ( .A(n648), .B(KEYINPUT87), .ZN(n649) );
  NOR2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n651), .A2(G48), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(G305) );
  XOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT90), .Z(n654) );
  XNOR2_X1 U740 ( .A(G288), .B(n654), .ZN(n655) );
  XNOR2_X1 U741 ( .A(G166), .B(n655), .ZN(n658) );
  XOR2_X1 U742 ( .A(n663), .B(G290), .Z(n656) );
  XNOR2_X1 U743 ( .A(n656), .B(G299), .ZN(n657) );
  XNOR2_X1 U744 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U745 ( .A(n659), .B(n955), .ZN(n660) );
  XNOR2_X1 U746 ( .A(n660), .B(G305), .ZN(n895) );
  XNOR2_X1 U747 ( .A(n661), .B(n895), .ZN(n662) );
  NAND2_X1 U748 ( .A1(n662), .A2(G868), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U759 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G96), .A2(n673), .ZN(n830) );
  NAND2_X1 U761 ( .A1(n830), .A2(G2106), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U764 ( .A1(G108), .A2(n675), .ZN(n831) );
  NAND2_X1 U765 ( .A1(n831), .A2(G567), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n832) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U768 ( .A1(n832), .A2(n678), .ZN(n679) );
  XOR2_X1 U769 ( .A(KEYINPUT91), .B(n679), .Z(n829) );
  NAND2_X1 U770 ( .A1(n829), .A2(G36), .ZN(G176) );
  INV_X1 U771 ( .A(n740), .ZN(n683) );
  NAND2_X1 U772 ( .A1(G1348), .A2(n722), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G2067), .A2(n708), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n691) );
  NOR2_X1 U775 ( .A1(n692), .A2(n691), .ZN(n690) );
  AND2_X1 U776 ( .A1(n708), .A2(G1996), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(KEYINPUT26), .ZN(n687) );
  NOR2_X1 U778 ( .A1(n688), .A2(n955), .ZN(n689) );
  NOR2_X1 U779 ( .A1(n690), .A2(n689), .ZN(n694) );
  AND2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n708), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n722), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U785 ( .A1(G299), .A2(n702), .ZN(n699) );
  XNOR2_X1 U786 ( .A(n699), .B(KEYINPUT98), .ZN(n700) );
  NOR2_X1 U787 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n702), .A2(G299), .ZN(n703) );
  XOR2_X1 U789 ( .A(KEYINPUT28), .B(n703), .Z(n704) );
  XNOR2_X1 U790 ( .A(n706), .B(KEYINPUT29), .ZN(n712) );
  NOR2_X1 U791 ( .A1(n708), .A2(G1961), .ZN(n707) );
  XNOR2_X1 U792 ( .A(n707), .B(KEYINPUT97), .ZN(n710) );
  XNOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .ZN(n977) );
  NAND2_X1 U794 ( .A1(n708), .A2(n977), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U796 ( .A1(G171), .A2(n714), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U798 ( .A1(G171), .A2(n714), .ZN(n715) );
  XNOR2_X1 U799 ( .A(n715), .B(KEYINPUT100), .ZN(n720) );
  NAND2_X1 U800 ( .A1(G8), .A2(n722), .ZN(n811) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n811), .ZN(n735) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n722), .ZN(n732) );
  NOR2_X1 U803 ( .A1(n735), .A2(n732), .ZN(n716) );
  NAND2_X1 U804 ( .A1(G8), .A2(n716), .ZN(n717) );
  XNOR2_X1 U805 ( .A(KEYINPUT30), .B(n717), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n718), .A2(G168), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n733), .A2(G286), .ZN(n727) );
  NOR2_X1 U809 ( .A1(G1971), .A2(n811), .ZN(n724) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n722), .ZN(n723) );
  NOR2_X1 U811 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U812 ( .A1(n725), .A2(G303), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U814 ( .A(KEYINPUT101), .B(n728), .Z(n729) );
  NAND2_X1 U815 ( .A1(n729), .A2(G8), .ZN(n731) );
  XNOR2_X1 U816 ( .A(n731), .B(n730), .ZN(n800) );
  NAND2_X1 U817 ( .A1(n732), .A2(G8), .ZN(n737) );
  INV_X1 U818 ( .A(n733), .ZN(n734) );
  NOR2_X1 U819 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U820 ( .A1(n737), .A2(n736), .ZN(n801) );
  NOR2_X1 U821 ( .A1(G1981), .A2(G305), .ZN(n738) );
  XOR2_X1 U822 ( .A(n738), .B(KEYINPUT24), .Z(n739) );
  NOR2_X1 U823 ( .A1(n811), .A2(n739), .ZN(n779) );
  NOR2_X1 U824 ( .A1(n779), .A2(n811), .ZN(n773) );
  NOR2_X1 U825 ( .A1(n741), .A2(n740), .ZN(n796) );
  XNOR2_X1 U826 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  XNOR2_X1 U827 ( .A(n742), .B(KEYINPUT92), .ZN(n794) );
  NAND2_X1 U828 ( .A1(G140), .A2(n875), .ZN(n744) );
  NAND2_X1 U829 ( .A1(G104), .A2(n876), .ZN(n743) );
  NAND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U831 ( .A(KEYINPUT34), .B(n745), .ZN(n752) );
  XNOR2_X1 U832 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n750) );
  NAND2_X1 U833 ( .A1(n870), .A2(G128), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n871), .A2(G116), .ZN(n746) );
  XOR2_X1 U835 ( .A(KEYINPUT93), .B(n746), .Z(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U837 ( .A(n750), .B(n749), .Z(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U839 ( .A(KEYINPUT36), .B(n753), .ZN(n892) );
  NOR2_X1 U840 ( .A1(n794), .A2(n892), .ZN(n1000) );
  NAND2_X1 U841 ( .A1(n796), .A2(n1000), .ZN(n791) );
  NAND2_X1 U842 ( .A1(n875), .A2(G131), .ZN(n756) );
  NAND2_X1 U843 ( .A1(G95), .A2(n876), .ZN(n754) );
  XOR2_X1 U844 ( .A(KEYINPUT95), .B(n754), .Z(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U846 ( .A1(G119), .A2(n870), .ZN(n758) );
  NAND2_X1 U847 ( .A1(G107), .A2(n871), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  OR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n885) );
  AND2_X1 U850 ( .A1(n885), .A2(G1991), .ZN(n770) );
  NAND2_X1 U851 ( .A1(G129), .A2(n870), .ZN(n761) );
  XNOR2_X1 U852 ( .A(n761), .B(KEYINPUT96), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G141), .A2(n875), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G117), .A2(n871), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n876), .A2(G105), .ZN(n764) );
  XOR2_X1 U857 ( .A(KEYINPUT38), .B(n764), .Z(n765) );
  NOR2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n867) );
  AND2_X1 U860 ( .A1(n867), .A2(G1996), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n1002) );
  INV_X1 U862 ( .A(n796), .ZN(n771) );
  NOR2_X1 U863 ( .A1(n1002), .A2(n771), .ZN(n788) );
  INV_X1 U864 ( .A(n788), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n791), .A2(n772), .ZN(n814) );
  NOR2_X1 U866 ( .A1(n773), .A2(n814), .ZN(n774) );
  XNOR2_X1 U867 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U868 ( .A1(n962), .A2(n796), .ZN(n818) );
  AND2_X1 U869 ( .A1(n774), .A2(n818), .ZN(n776) );
  AND2_X1 U870 ( .A1(n801), .A2(n776), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n800), .A2(n775), .ZN(n785) );
  INV_X1 U872 ( .A(n776), .ZN(n783) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U874 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U875 ( .A(n778), .B(KEYINPUT104), .ZN(n781) );
  INV_X1 U876 ( .A(n779), .ZN(n780) );
  AND2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n799) );
  NOR2_X1 U880 ( .A1(G1996), .A2(n867), .ZN(n1008) );
  NOR2_X1 U881 ( .A1(G1986), .A2(G290), .ZN(n786) );
  NOR2_X1 U882 ( .A1(G1991), .A2(n885), .ZN(n996) );
  NOR2_X1 U883 ( .A1(n786), .A2(n996), .ZN(n787) );
  NOR2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U885 ( .A1(n1008), .A2(n789), .ZN(n790) );
  XNOR2_X1 U886 ( .A(n790), .B(KEYINPUT39), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U888 ( .A(KEYINPUT105), .B(n793), .Z(n795) );
  NAND2_X1 U889 ( .A1(n794), .A2(n892), .ZN(n1012) );
  NAND2_X1 U890 ( .A1(n795), .A2(n1012), .ZN(n797) );
  AND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n824) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n805) );
  NOR2_X1 U894 ( .A1(G1976), .A2(G288), .ZN(n809) );
  NOR2_X1 U895 ( .A1(G1971), .A2(G303), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n809), .A2(n802), .ZN(n947) );
  INV_X1 U897 ( .A(KEYINPUT33), .ZN(n803) );
  AND2_X1 U898 ( .A1(n947), .A2(n803), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n822) );
  NAND2_X1 U900 ( .A1(G288), .A2(G1976), .ZN(n806) );
  XOR2_X1 U901 ( .A(KEYINPUT103), .B(n806), .Z(n946) );
  INV_X1 U902 ( .A(n946), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n807), .A2(n811), .ZN(n808) );
  NOR2_X1 U904 ( .A1(KEYINPUT33), .A2(n808), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n809), .A2(KEYINPUT33), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n817) );
  XOR2_X1 U908 ( .A(G1981), .B(G305), .Z(n943) );
  INV_X1 U909 ( .A(n814), .ZN(n815) );
  AND2_X1 U910 ( .A1(n943), .A2(n815), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n820) );
  INV_X1 U912 ( .A(n818), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U916 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U919 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(G188) );
  XOR2_X1 U922 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n832), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT109), .B(G2678), .Z(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2090), .Z(n836) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2096), .B(G2100), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U938 ( .A(G2078), .B(G2084), .Z(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1976), .B(G1956), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1991), .B(G1961), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT41), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(n851), .ZN(n852) );
  XOR2_X1 U950 ( .A(n852), .B(G1996), .Z(G229) );
  NAND2_X1 U951 ( .A1(G136), .A2(n875), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G112), .A2(n871), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U954 ( .A1(n870), .A2(G124), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G100), .A2(n876), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G130), .A2(n870), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G118), .A2(n871), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G142), .A2(n875), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G106), .A2(n876), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n864), .B(KEYINPUT45), .Z(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n869), .B(n995), .Z(n884) );
  NAND2_X1 U969 ( .A1(G127), .A2(n870), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G115), .A2(n871), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U973 ( .A1(G139), .A2(n875), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G103), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(KEYINPUT112), .B(n879), .Z(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n882), .B(KEYINPUT113), .ZN(n1003) );
  XNOR2_X1 U979 ( .A(n1003), .B(G162), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n889) );
  XOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n887) );
  XOR2_X1 U982 ( .A(n885), .B(KEYINPUT46), .Z(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(n889), .B(n888), .Z(n891) );
  XNOR2_X1 U985 ( .A(G164), .B(G160), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U989 ( .A(n895), .B(n958), .Z(n897) );
  XNOR2_X1 U990 ( .A(G286), .B(G171), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  XNOR2_X1 U993 ( .A(G2451), .B(G2443), .ZN(n908) );
  XOR2_X1 U994 ( .A(G2446), .B(G2454), .Z(n900) );
  XNOR2_X1 U995 ( .A(KEYINPUT106), .B(G2435), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U997 ( .A(KEYINPUT107), .B(G2438), .Z(n902) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G2430), .B(G2427), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n909), .A2(G14), .ZN(n915) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n915), .ZN(G401) );
  XOR2_X1 U1014 ( .A(G16), .B(KEYINPUT122), .Z(n940) );
  XOR2_X1 U1015 ( .A(G1986), .B(G24), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G1971), .B(G22), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G23), .B(G1976), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1961), .B(G5), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G21), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(G1341), .B(G19), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(G1981), .B(G6), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1029 ( .A(KEYINPUT123), .B(n928), .Z(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n929), .B(G4), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n930), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(G20), .B(G1956), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT60), .B(n935), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT61), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT126), .ZN(n968) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(KEYINPUT120), .ZN(n966) );
  XNOR2_X1 U1043 ( .A(G168), .B(G1966), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT57), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(G303), .A2(G1971), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G299), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n952), .B(KEYINPUT121), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n958), .B(G1348), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G171), .B(G1961), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT127), .B(n969), .ZN(n994) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n970), .ZN(n988) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n986) );
  XNOR2_X1 U1066 ( .A(KEYINPUT115), .B(G2067), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n971), .B(G26), .ZN(n976) );
  XOR2_X1 U1068 ( .A(G25), .B(G1991), .Z(n972) );
  NAND2_X1 U1069 ( .A1(n972), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n982) );
  XOR2_X1 U1073 ( .A(n977), .B(G27), .Z(n979) );
  XNOR2_X1 U1074 ( .A(G1996), .B(G32), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1076 ( .A(n980), .B(KEYINPUT116), .Z(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1078 ( .A(KEYINPUT53), .B(n983), .Z(n984) );
  XNOR2_X1 U1079 ( .A(n984), .B(KEYINPUT117), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT118), .ZN(n990) );
  XOR2_X1 U1083 ( .A(KEYINPUT55), .B(n990), .Z(n992) );
  XNOR2_X1 U1084 ( .A(G29), .B(KEYINPUT119), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1021) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1015) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1003), .Z(n1005) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1006), .Z(n1011) );
  XOR2_X1 U1096 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .Z(n1017) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1017), .ZN(n1019) );
  INV_X1 U1104 ( .A(G29), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(G11), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

