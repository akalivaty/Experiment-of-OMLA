//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n204), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(new_n233));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OR2_X1    g0046(.A1(KEYINPUT70), .A2(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT70), .A2(G1), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n247), .A2(G13), .A3(G20), .A4(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT70), .A2(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT70), .A2(G1), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n250), .A2(new_n251), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n254), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n210), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G159), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT78), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT78), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(G159), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G58), .ZN(new_n271));
  INV_X1    g0071(.A(G68), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n273), .B2(new_n203), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT77), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n283), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n276), .A2(new_n210), .A3(new_n277), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT7), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n275), .B1(new_n288), .B2(G68), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n262), .B1(new_n289), .B2(KEYINPUT16), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT16), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n272), .B1(new_n287), .B2(new_n278), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n261), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n263), .C2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(G226), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT79), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(new_n277), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n301), .A2(KEYINPUT79), .A3(G226), .A4(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(G223), .B(new_n304), .C1(new_n281), .C2(new_n282), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n297), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n247), .A2(new_n248), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G41), .A2(G45), .ZN(new_n311));
  OAI211_X1 g0111(.A(G232), .B(new_n297), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G1), .ZN(new_n314));
  OR2_X1    g0114(.A1(KEYINPUT69), .A2(G41), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT69), .A2(G41), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(G45), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n295), .B1(new_n309), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT80), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT80), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n312), .A2(new_n322), .A3(new_n318), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n307), .B1(new_n300), .B2(new_n302), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n323), .C1(new_n297), .C2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT71), .B(G179), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n294), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT18), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n309), .B2(new_n319), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n325), .B2(G190), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n294), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n253), .B1(G33), .B2(G41), .ZN(new_n337));
  INV_X1    g0137(.A(new_n311), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n258), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G226), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(new_n318), .ZN(new_n341));
  AOI21_X1  g0141(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G222), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n301), .A2(G223), .A3(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G77), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n301), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT72), .B1(new_n349), .B2(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n326), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n249), .A2(new_n262), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(G50), .A3(new_n259), .ZN(new_n355));
  INV_X1    g0155(.A(G50), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n250), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n210), .A2(G33), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n251), .A2(new_n358), .B1(new_n359), .B2(new_n264), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n254), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT72), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n352), .B(new_n363), .C1(new_n364), .C2(new_n351), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n310), .A2(new_n210), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n353), .A2(new_n366), .A3(new_n345), .ZN(new_n367));
  INV_X1    g0167(.A(new_n251), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n371), .B2(new_n254), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n249), .A2(G77), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n301), .A2(G232), .A3(new_n304), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n301), .A2(G238), .A3(G1698), .ZN(new_n378));
  INV_X1    g0178(.A(G107), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n301), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n337), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n339), .A2(G244), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n318), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G200), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n376), .B(new_n384), .C1(new_n385), .C2(new_n383), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n383), .A2(new_n327), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n295), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n375), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n363), .A2(KEYINPUT9), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n363), .A2(KEYINPUT9), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(G200), .B2(new_n348), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT10), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n348), .B2(new_n385), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n341), .A2(new_n347), .A3(KEYINPUT74), .A4(G190), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n393), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n394), .B1(new_n393), .B2(new_n398), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n365), .B(new_n390), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n354), .A2(G68), .A3(new_n259), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n272), .A2(G20), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n404), .B1(new_n358), .B2(new_n345), .C1(new_n356), .C2(new_n264), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n254), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(KEYINPUT11), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT11), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n405), .B2(new_n254), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n249), .A2(G68), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n402), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n406), .B(KEYINPUT11), .ZN(new_n414));
  INV_X1    g0214(.A(new_n412), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT76), .A4(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n342), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n301), .A2(G232), .A3(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n297), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(G238), .B(new_n297), .C1(new_n310), .C2(new_n311), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n318), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT13), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n342), .A2(G226), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n420), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n337), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  INV_X1    g0229(.A(new_n423), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(G169), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n424), .A2(new_n431), .A3(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n432), .B2(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n418), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(G200), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n410), .A2(new_n412), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n385), .C2(new_n432), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n336), .A2(new_n401), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT83), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT5), .B1(new_n315), .B2(new_n316), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n247), .A2(G45), .A3(new_n248), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n256), .A2(new_n257), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT69), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT69), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n451), .A2(G41), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n337), .A2(new_n313), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n456), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G257), .A3(new_n297), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  OAI211_X1 g0263(.A(G250), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n464));
  OAI211_X1 g0264(.A(G244), .B(new_n304), .C1(new_n281), .C2(new_n282), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT4), .B1(new_n342), .B2(G244), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n337), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT85), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n458), .A4(new_n461), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G190), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n249), .A2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n247), .A2(G33), .A3(new_n248), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n354), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n480), .A2(G97), .A3(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n379), .A2(KEYINPUT81), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n379), .A2(KEYINPUT81), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT81), .B(G107), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(G97), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n490), .A3(G20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n267), .A2(G77), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT82), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n287), .A2(new_n278), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n479), .B1(new_n498), .B2(new_n254), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n458), .A2(new_n500), .A3(new_n461), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n458), .B2(new_n461), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n469), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n473), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n496), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n254), .B1(new_n506), .B2(new_n493), .ZN(new_n507));
  INV_X1    g0307(.A(new_n479), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  INV_X1    g0310(.A(new_n467), .ZN(new_n511));
  INV_X1    g0311(.A(new_n468), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n297), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n458), .A2(new_n461), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n295), .A3(new_n471), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n326), .B(new_n469), .C1(new_n501), .C2(new_n502), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n509), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n505), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n249), .A2(G107), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n520), .A2(KEYINPUT25), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n379), .B2(new_n477), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n301), .A2(new_n210), .A3(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT22), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n301), .A2(new_n527), .A3(new_n210), .A4(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n358), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n210), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n379), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT24), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n524), .B1(new_n540), .B2(new_n254), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT95), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n460), .A2(G264), .A3(new_n297), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(new_n304), .C1(new_n281), .C2(new_n282), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G294), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n337), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n543), .A2(new_n548), .A3(KEYINPUT93), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT93), .B1(new_n543), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(G200), .B1(new_n551), .B2(new_n458), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n458), .A2(new_n543), .A3(new_n548), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n541), .B(new_n542), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n543), .A2(new_n548), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n543), .A2(new_n548), .A3(KEYINPUT93), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n458), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n554), .B1(new_n560), .B2(new_n331), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n529), .A2(new_n538), .A3(new_n535), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n538), .B1(new_n529), .B2(new_n535), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n254), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n477), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT95), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n210), .B(G68), .C1(new_n281), .C2(new_n282), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n358), .B2(new_n478), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g0374(.A1(KEYINPUT87), .A2(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(KEYINPUT87), .A2(G87), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n487), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n210), .B1(new_n426), .B2(new_n572), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n262), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n370), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n249), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n570), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n571), .A3(new_n573), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(new_n254), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n583), .A2(new_n586), .B1(new_n581), .B2(new_n565), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n247), .A2(G45), .A3(new_n313), .A4(new_n248), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n297), .B(new_n589), .C1(new_n450), .C2(G250), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT86), .ZN(new_n591));
  INV_X1    g0391(.A(G250), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n337), .B1(new_n447), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n342), .A2(G238), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n301), .A2(G244), .A3(G1698), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n337), .ZN(new_n601));
  AOI21_X1  g0401(.A(G169), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n591), .A2(new_n595), .B1(new_n600), .B2(new_n337), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n326), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n596), .A2(G190), .A3(new_n601), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n331), .B1(new_n596), .B2(new_n601), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n249), .A2(new_n262), .A3(new_n476), .A4(G87), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT89), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n583), .B2(new_n586), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n588), .A2(new_n604), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n519), .A2(new_n569), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n558), .A2(G179), .A3(new_n458), .A4(new_n559), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n553), .A2(G169), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(KEYINPUT94), .A3(new_n614), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n567), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n460), .A2(G270), .A3(new_n297), .ZN(new_n621));
  OAI211_X1 g0421(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n622));
  OAI211_X1 g0422(.A(G257), .B(new_n304), .C1(new_n281), .C2(new_n282), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n337), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n458), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n250), .A2(new_n530), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n249), .A2(new_n262), .A3(new_n476), .A4(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n463), .B(new_n210), .C1(G33), .C2(new_n478), .ZN(new_n632));
  AOI221_X4 g0432(.A(KEYINPUT90), .B1(new_n530), .B2(G20), .C1(new_n252), .C2(new_n253), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n530), .A2(G20), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n254), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(KEYINPUT20), .B(new_n632), .C1(new_n633), .C2(new_n636), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n620), .B1(new_n628), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT92), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT92), .B(new_n620), .C1(new_n628), .C2(new_n641), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n627), .A2(KEYINPUT21), .A3(G169), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n458), .A2(new_n621), .A3(new_n626), .A4(G179), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n627), .A2(new_n385), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n627), .A2(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n641), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n649), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n619), .A2(new_n650), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n444), .A2(new_n612), .A3(new_n656), .ZN(G372));
  INV_X1    g0457(.A(new_n365), .ZN(new_n658));
  INV_X1    g0458(.A(new_n438), .ZN(new_n659));
  INV_X1    g0459(.A(new_n389), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n441), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n335), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n330), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n399), .A2(new_n400), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n631), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n254), .A2(new_n635), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n254), .A2(new_n634), .A3(new_n635), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT20), .B1(new_n670), .B2(new_n632), .ZN(new_n671));
  INV_X1    g0471(.A(new_n640), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(G169), .A3(new_n627), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT92), .B1(new_n674), .B2(new_n620), .ZN(new_n675));
  INV_X1    g0475(.A(new_n645), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n654), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT96), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT96), .B(new_n654), .C1(new_n675), .C2(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n567), .A2(new_n615), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n519), .A2(new_n569), .A3(new_n611), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n679), .A2(KEYINPUT97), .A3(new_n680), .A4(new_n681), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n596), .A2(new_n326), .A3(new_n601), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n603), .B2(G169), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n587), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n509), .A2(new_n516), .A3(new_n517), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n611), .A2(new_n691), .A3(KEYINPUT26), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n583), .A2(new_n586), .ZN(new_n694));
  INV_X1    g0494(.A(new_n609), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n596), .A2(G190), .A3(new_n601), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n603), .B2(new_n331), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n696), .A2(new_n698), .B1(new_n689), .B2(new_n587), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n693), .B1(new_n699), .B2(new_n518), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n690), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n665), .B1(new_n703), .B2(new_n444), .ZN(G369));
  AND2_X1   g0504(.A1(new_n210), .A2(G13), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n258), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G213), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G343), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n679), .A2(new_n673), .A3(new_n680), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n650), .A2(new_n655), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n673), .A2(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n712), .A2(new_n653), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n711), .B1(new_n617), .B2(new_n618), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n569), .B1(new_n541), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n711), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n619), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n713), .A2(new_n720), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n567), .A2(new_n615), .A3(new_n720), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n723), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n213), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n317), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n577), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n217), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n734), .A2(KEYINPUT98), .B1(new_n735), .B2(new_n730), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(KEYINPUT98), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n702), .A2(new_n720), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n619), .A2(new_n650), .A3(new_n655), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n701), .B1(new_n612), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .A3(new_n720), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n656), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n685), .A2(new_n746), .A3(new_n720), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n470), .A2(new_n472), .ZN(new_n749));
  INV_X1    g0549(.A(new_n648), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n551), .A2(new_n603), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n515), .A2(new_n471), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n596), .A2(new_n601), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n648), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT30), .A4(new_n551), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n627), .A2(new_n326), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT99), .B2(new_n754), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(new_n560), .A4(new_n503), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n752), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n761), .B2(new_n711), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G330), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT100), .B1(new_n745), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT100), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n741), .C2(new_n744), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n738), .B1(new_n773), .B2(G1), .ZN(G364));
  INV_X1    g0574(.A(new_n717), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n209), .B1(new_n705), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n730), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT101), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n717), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n716), .A2(G330), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n776), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n253), .B1(G20), .B2(new_n295), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n385), .A2(G179), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n210), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n326), .A2(new_n210), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n790), .B1(new_n794), .B2(new_n272), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT103), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n385), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(G179), .B1(new_n797), .B2(KEYINPUT102), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(KEYINPUT102), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G159), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT32), .Z(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(new_n331), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n379), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n210), .A2(new_n385), .A3(new_n331), .A4(G179), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n575), .A2(new_n576), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n283), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n385), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n791), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G190), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n791), .A2(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n808), .B1(new_n810), .B2(new_n271), .C1(new_n345), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n792), .A2(new_n385), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n805), .B(new_n813), .C1(G50), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n796), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n301), .B1(new_n806), .B2(G303), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n788), .C1(new_n812), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n810), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G322), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n793), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n803), .A2(G283), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n814), .A2(G326), .B1(new_n800), .B2(G329), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n786), .B1(new_n816), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n785), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n213), .A2(new_n283), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n449), .B2(new_n735), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n245), .B2(new_n449), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n213), .A2(new_n301), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(G116), .B2(new_n213), .C1(new_n207), .C2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n780), .B(new_n828), .C1(new_n832), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT104), .ZN(new_n839));
  INV_X1    g0639(.A(new_n831), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n716), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n784), .A2(new_n841), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n785), .A2(new_n829), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n375), .A2(new_n711), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n386), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n389), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n660), .A2(new_n720), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n779), .B1(G77), .B2(new_n844), .C1(new_n849), .C2(new_n830), .ZN(new_n850));
  INV_X1    g0650(.A(new_n812), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n821), .B1(new_n851), .B2(G159), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G137), .A2(new_n814), .B1(new_n793), .B2(G150), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(KEYINPUT105), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(KEYINPUT105), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  INV_X1    g0659(.A(new_n806), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n301), .B1(new_n271), .B2(new_n788), .C1(new_n860), .C2(new_n356), .ZN(new_n861));
  INV_X1    g0661(.A(new_n800), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n861), .B(new_n864), .C1(G68), .C2(new_n803), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n803), .A2(G87), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G283), .B2(new_n793), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n301), .B1(new_n806), .B2(G107), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n790), .B(new_n869), .C1(new_n530), .C2(new_n812), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(G294), .B2(new_n821), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n814), .A2(G303), .B1(new_n800), .B2(G311), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n786), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n850), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n847), .A2(new_n848), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n739), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n390), .A2(new_n720), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n687), .B2(new_n701), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n779), .B1(new_n881), .B2(new_n767), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(new_n770), .A3(new_n880), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  NOR2_X1   g0685(.A1(new_n216), .A2(new_n530), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n485), .A2(new_n490), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT35), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  OR3_X1    g0691(.A1(new_n217), .A2(new_n345), .A3(new_n273), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n201), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(G13), .B(new_n258), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n288), .A2(G68), .ZN(new_n897));
  INV_X1    g0697(.A(new_n275), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(KEYINPUT16), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n293), .A3(new_n254), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n333), .A2(new_n900), .A3(new_n260), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n329), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT107), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n294), .B2(new_n709), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n260), .ZN(new_n905));
  INV_X1    g0705(.A(new_n709), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT107), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT107), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n903), .B(new_n709), .C1(new_n900), .C2(new_n260), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n322), .B1(new_n312), .B2(new_n318), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n312), .A2(new_n322), .A3(new_n318), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n309), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n318), .B(new_n312), .C1(new_n324), .C2(new_n297), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n916), .A2(new_n326), .B1(new_n295), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n334), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT108), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n913), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n919), .A2(new_n920), .A3(new_n334), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT108), .B1(new_n924), .B2(new_n908), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n910), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n908), .B1(new_n330), .B2(new_n335), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n290), .B1(KEYINPUT16), .B2(new_n289), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n260), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n906), .B1(new_n294), .B2(new_n333), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n918), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n922), .B1(new_n913), .B2(new_n921), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT108), .A4(new_n920), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n931), .A2(new_n906), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n330), .B2(new_n335), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n896), .B1(new_n929), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n659), .A2(new_n720), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n934), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n923), .B2(new_n925), .ZN(new_n946));
  INV_X1    g0746(.A(new_n940), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT38), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n938), .B1(new_n937), .B2(new_n940), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT39), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n949), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n418), .A2(new_n711), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n438), .A2(new_n441), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n438), .B2(new_n441), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n848), .B(KEYINPUT106), .Z(new_n958));
  OAI211_X1 g0758(.A(new_n952), .B(new_n957), .C1(new_n879), .C2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n330), .A2(new_n906), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n951), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n711), .B1(new_n687), .B2(new_n701), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n744), .B(new_n443), .C1(new_n962), .C2(KEYINPUT29), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n665), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n961), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n849), .B1(new_n954), .B2(new_n955), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n747), .B2(new_n765), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n952), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  INV_X1    g0769(.A(new_n955), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n438), .A2(new_n441), .A3(new_n953), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n876), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n612), .A2(new_n656), .A3(new_n711), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n761), .A2(new_n711), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT31), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n762), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n972), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n969), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n935), .A2(new_n936), .B1(KEYINPUT37), .B2(new_n909), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n938), .B1(new_n980), .B2(new_n927), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n948), .A2(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n968), .A2(new_n969), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n973), .A2(new_n977), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n444), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n443), .A3(new_n766), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(G330), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n965), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n258), .B2(new_n705), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n965), .A2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n895), .B1(new_n990), .B2(new_n991), .ZN(G367));
  INV_X1    g0792(.A(new_n232), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n832), .B1(new_n213), .B2(new_n370), .C1(new_n993), .C2(new_n833), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n779), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n814), .A2(G143), .B1(new_n800), .B2(G137), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n345), .B2(new_n804), .C1(new_n265), .C2(new_n794), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n789), .A2(G68), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n283), .B1(new_n806), .B2(G58), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n359), .B2(new_n810), .C1(new_n201), .C2(new_n812), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n860), .B2(new_n530), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n283), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G107), .B2(new_n789), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G283), .A2(new_n851), .B1(new_n821), .B2(G303), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G294), .A2(new_n793), .B1(new_n814), .B2(G311), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n806), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT110), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n800), .A2(G317), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n803), .A2(G97), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n997), .A2(new_n1001), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n995), .B1(new_n1015), .B2(new_n785), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n696), .A2(new_n711), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1017), .A2(new_n587), .A3(new_n689), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n611), .B2(new_n1017), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n831), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n519), .B1(new_n499), .B2(new_n720), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n691), .A2(new_n711), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(new_n725), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n518), .B1(new_n1022), .B2(new_n619), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n720), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(KEYINPUT109), .B1(KEYINPUT42), .B2(new_n1026), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1030), .A2(KEYINPUT109), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT43), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1031), .A2(new_n1032), .B1(new_n1033), .B2(new_n1019), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1019), .A2(new_n1033), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n723), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n1025), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1036), .B(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n727), .A2(new_n1025), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT44), .Z(new_n1041));
  NOR2_X1   g0841(.A1(new_n727), .A2(new_n1025), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT45), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1037), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1041), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n722), .A2(new_n724), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n725), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n776), .A2(new_n782), .A3(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n717), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n773), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n730), .B(KEYINPUT41), .Z(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n778), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1021), .B1(new_n1039), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT112), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(G387));
  NAND2_X1  g0859(.A1(new_n745), .A2(new_n767), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n769), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n745), .A2(KEYINPUT100), .A3(new_n767), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n1062), .A3(new_n1052), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1052), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n768), .B2(new_n771), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1065), .A3(new_n730), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n722), .A2(new_n831), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n237), .A2(new_n449), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1068), .A2(new_n833), .B1(new_n732), .B2(new_n836), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n251), .A2(G50), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n732), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1069), .A2(new_n1074), .B1(new_n379), .B2(new_n729), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n832), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n779), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n793), .A2(new_n368), .B1(new_n851), .B2(G68), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT114), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n821), .A2(G50), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n789), .A2(new_n581), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n283), .B1(new_n806), .B2(G77), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n1012), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n814), .A2(G159), .B1(new_n800), .B2(G150), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1079), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n301), .B1(new_n800), .B2(G326), .ZN(new_n1086));
  INV_X1    g0886(.A(G283), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n860), .A2(new_n818), .B1(new_n1087), .B2(new_n788), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G303), .A2(new_n851), .B1(new_n821), .B2(G317), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n814), .A2(G322), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n819), .C2(new_n794), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1086), .B1(new_n530), .B2(new_n804), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1085), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1077), .B1(new_n1098), .B2(new_n785), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1064), .A2(new_n778), .B1(new_n1067), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1066), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT115), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT115), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1066), .A2(new_n1103), .A3(new_n1100), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(G393));
  INV_X1    g0905(.A(new_n1065), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1046), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n1044), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n731), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT116), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n777), .B1(new_n1047), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1111), .B2(new_n1047), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n814), .A2(G317), .B1(new_n821), .B2(G311), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  OAI221_X1 g0915(.A(new_n283), .B1(new_n530), .B2(new_n788), .C1(new_n860), .C2(new_n1087), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1116), .B(new_n805), .C1(G294), .C2(new_n851), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n793), .A2(G303), .B1(new_n800), .B2(G322), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n814), .A2(G150), .B1(new_n821), .B2(G159), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT51), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n789), .A2(G77), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n301), .C1(new_n272), .C2(new_n860), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1123), .B(new_n867), .C1(new_n368), .C2(new_n851), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n793), .A2(new_n202), .B1(new_n800), .B2(G143), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n786), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n242), .A2(new_n833), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1076), .B1(G97), .B2(new_n729), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n780), .B(new_n1127), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1024), .B2(new_n840), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1110), .A2(new_n1113), .A3(new_n1131), .ZN(G390));
  NOR3_X1   g0932(.A1(new_n767), .A2(new_n876), .A3(new_n956), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n943), .B1(new_n929), .B2(new_n941), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n743), .A2(new_n720), .A3(new_n849), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n958), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n956), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n944), .B1(new_n948), .B2(new_n981), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n611), .A2(new_n518), .A3(new_n505), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n619), .A2(new_n650), .A3(new_n655), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n569), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n711), .B(new_n876), .C1(new_n1143), .C2(new_n701), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n957), .B1(new_n1144), .B2(new_n958), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT117), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n957), .B1(new_n879), .B2(new_n958), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n943), .B1(new_n942), .B2(new_n950), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1133), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n943), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n942), .A2(new_n950), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1138), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1140), .A2(new_n1145), .A3(KEYINPUT117), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1133), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n443), .B(G330), .C1(new_n973), .C2(new_n977), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n766), .A2(KEYINPUT118), .A3(G330), .A4(new_n443), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n963), .A3(new_n665), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n880), .A2(new_n1136), .ZN(new_n1166));
  INV_X1    g0966(.A(G330), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n985), .A2(new_n1167), .A3(new_n876), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n957), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1169), .B2(new_n1133), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1168), .B2(new_n957), .ZN(new_n1172));
  OAI211_X1 g0972(.A(KEYINPUT119), .B(G330), .C1(new_n973), .C2(new_n977), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n849), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT119), .B1(new_n766), .B2(G330), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n956), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1165), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1159), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1150), .A2(new_n1158), .A3(new_n1178), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n730), .A3(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1152), .A2(new_n829), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n779), .B1(new_n368), .B2(new_n844), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n301), .B1(new_n806), .B2(G87), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1122), .B(new_n1186), .C1(new_n530), .C2(new_n810), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G97), .B2(new_n851), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G68), .A2(new_n803), .B1(new_n800), .B2(G294), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G107), .A2(new_n793), .B1(new_n814), .B2(G283), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n806), .A2(G150), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT53), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n301), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G132), .B2(new_n821), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n814), .A2(G128), .B1(new_n800), .B2(G125), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n201), .C2(new_n804), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT54), .B(G143), .Z(new_n1198));
  AOI22_X1  g0998(.A1(new_n851), .A2(new_n1198), .B1(G159), .B2(new_n789), .ZN(new_n1199));
  INV_X1    g0999(.A(G137), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n794), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1191), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1185), .B1(new_n1203), .B2(new_n785), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1183), .A2(new_n778), .B1(new_n1184), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1182), .A2(new_n1205), .ZN(G378));
  INV_X1    g1006(.A(new_n1165), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n951), .A2(new_n959), .A3(new_n960), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n664), .A2(new_n365), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n363), .A2(new_n906), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n983), .B2(G330), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n967), .B(KEYINPUT40), .C1(new_n929), .C2(new_n941), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n978), .B1(new_n948), .B2(new_n949), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(G330), .C1(new_n1223), .C2(KEYINPUT40), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1210), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n983), .A2(new_n1220), .A3(G330), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n961), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1209), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1208), .A2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1181), .A2(new_n1207), .B1(new_n1230), .B2(new_n1227), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n730), .C1(KEYINPUT57), .C2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1228), .A2(new_n961), .A3(new_n1229), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n961), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n778), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n780), .B1(new_n201), .B2(new_n843), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n851), .A2(G137), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n789), .A2(G150), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n806), .A2(new_n1198), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n814), .A2(G125), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n794), .B2(new_n863), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(G128), .C2(new_n821), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT121), .B(G124), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n263), .B(new_n296), .C1(new_n862), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G159), .B2(new_n803), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n821), .A2(G107), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n806), .A2(G77), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n301), .A2(new_n317), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n998), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n814), .A2(G116), .B1(new_n800), .B2(G283), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n803), .A2(G58), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n478), .C2(new_n794), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1256), .B(new_n1259), .C1(new_n581), .C2(new_n851), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT58), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1260), .A2(KEYINPUT58), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n356), .B1(G33), .B2(G41), .C1(new_n301), .C2(new_n317), .ZN(new_n1263));
  AND4_X1   g1063(.A1(new_n1252), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1238), .B1(new_n786), .B2(new_n1264), .C1(new_n1220), .C2(new_n830), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1237), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1234), .A2(new_n1267), .ZN(G375));
  NAND3_X1  g1068(.A1(new_n1170), .A2(new_n1177), .A3(new_n1165), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1179), .A2(new_n1055), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n956), .A2(new_n829), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n779), .B1(G68), .B2(new_n844), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT122), .Z(new_n1274));
  OAI221_X1 g1074(.A(new_n1081), .B1(new_n478), .B2(new_n860), .C1(new_n812), .C2(new_n379), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G283), .B2(new_n821), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n814), .A2(G294), .B1(new_n800), .B2(G303), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(new_n530), .C2(new_n794), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n301), .B1(new_n803), .B2(G77), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT123), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n301), .B1(new_n356), .B2(new_n788), .C1(new_n860), .C2(new_n265), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G137), .B2(new_n821), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n359), .B2(new_n812), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(G132), .A2(new_n814), .B1(new_n793), .B2(new_n1198), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n800), .A2(G128), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1258), .A3(new_n1285), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1278), .A2(new_n1280), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1274), .B1(new_n1287), .B2(new_n785), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1271), .A2(new_n778), .B1(new_n1272), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1270), .A2(new_n1289), .ZN(G381));
  XNOR2_X1  g1090(.A(G375), .B(KEYINPUT124), .ZN(new_n1291));
  INV_X1    g1091(.A(G396), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1102), .A2(new_n1292), .A3(new_n1104), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1270), .A2(new_n884), .A3(new_n1289), .ZN(new_n1294));
  NOR4_X1   g1094(.A1(G390), .A2(new_n1293), .A3(G378), .A4(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1058), .A2(new_n1291), .A3(new_n1295), .ZN(G407));
  INV_X1    g1096(.A(G378), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1291), .A2(G213), .A3(new_n710), .A4(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G407), .A2(G213), .A3(new_n1298), .ZN(G409));
  INV_X1    g1099(.A(new_n1057), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1104), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1103), .B1(new_n1066), .B2(new_n1100), .ZN(new_n1302));
  OAI21_X1  g1102(.A(G396), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1293), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT112), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G390), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1113), .A2(new_n1131), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1110), .A2(new_n1307), .B1(new_n1303), .B2(new_n1293), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1300), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(G390), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT112), .B1(new_n1303), .B2(new_n1293), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1310), .B(new_n1057), .C1(G390), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n710), .A2(G213), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1271), .A2(new_n1207), .A3(new_n1315), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1316), .A2(new_n729), .A3(new_n317), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1269), .B1(new_n1178), .B2(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1319), .B2(new_n1289), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1289), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n884), .B(new_n1321), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1234), .A2(G378), .A3(new_n1267), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1054), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1208), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1266), .B1(KEYINPUT125), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1208), .A2(new_n1325), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G378), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1314), .B(new_n1323), .C1(new_n1324), .C2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1234), .A2(G378), .A3(new_n1267), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1326), .A2(KEYINPUT125), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1335), .A2(new_n1267), .A3(new_n1329), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1334), .B1(new_n1336), .B2(G378), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1337), .A2(KEYINPUT62), .A3(new_n1314), .A4(new_n1323), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1333), .A2(KEYINPUT127), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1331), .A2(new_n1340), .A3(new_n1332), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n710), .A2(G213), .A3(G2897), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1320), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1319), .A2(G384), .A3(new_n1289), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1342), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1320), .A2(new_n1322), .A3(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1314), .B1(new_n1324), .B2(new_n1330), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1341), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1313), .B1(new_n1339), .B2(new_n1352), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1331), .A2(KEYINPUT63), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1331), .A2(KEYINPUT63), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1354), .B(new_n1355), .C1(new_n1356), .C2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1353), .A2(new_n1358), .ZN(G405));
  NAND2_X1  g1159(.A1(G375), .A2(new_n1297), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1334), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1361), .B(new_n1323), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1362), .B(new_n1313), .ZN(G402));
endmodule


