//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  XNOR2_X1  g000(.A(G134gat), .B(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G43gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT15), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT93), .B(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT94), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT94), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n209), .B2(new_n210), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n210), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n220), .B(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n208), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n214), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT96), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n207), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n205), .B(KEYINPUT97), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT15), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT95), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT95), .A4(KEYINPUT15), .ZN(new_n232));
  OR4_X1    g031(.A1(KEYINPUT98), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT98), .A3(new_n221), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n225), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT99), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n235), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n227), .A2(new_n228), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n215), .B(new_n238), .C1(KEYINPUT15), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n208), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n220), .B(new_n221), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n225), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  INV_X1    g047(.A(G92gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(KEYINPUT8), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT7), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n248), .B2(new_n249), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G99gat), .B(G106gat), .Z(new_n255));
  OR2_X1    g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT41), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n237), .A2(new_n264), .A3(new_n245), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT17), .B1(new_n224), .B2(new_n236), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n263), .A2(new_n267), .A3(KEYINPUT108), .ZN(new_n268));
  XNOR2_X1  g067(.A(G190gat), .B(G218gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT107), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT106), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n261), .A2(KEYINPUT41), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n267), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT108), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n246), .A2(new_n259), .B1(KEYINPUT41), .B2(new_n261), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT108), .B1(new_n263), .B2(new_n267), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n270), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n272), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n272), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n203), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n272), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n273), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(new_n274), .A3(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n202), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT16), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(G1gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT100), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n291), .B(new_n292), .C1(G1gat), .C2(new_n289), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(G8gat), .C1(new_n292), .C2(new_n291), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT101), .B1(new_n289), .B2(G1gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n291), .ZN(new_n296));
  INV_X1    g095(.A(G8gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT101), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(new_n265), .B2(new_n266), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n237), .B2(new_n245), .ZN(new_n303));
  NAND2_X1  g102(.A1(G229gat), .A2(G233gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT102), .Z(new_n305));
  NOR3_X1   g104(.A1(new_n301), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n246), .B(new_n300), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n305), .B(KEYINPUT13), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n306), .A2(KEYINPUT18), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT104), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT103), .B(KEYINPUT18), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n265), .A2(new_n266), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n302), .ZN(new_n316));
  INV_X1    g115(.A(new_n303), .ZN(new_n317));
  INV_X1    g116(.A(new_n305), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT104), .A3(new_n312), .ZN(new_n320));
  XOR2_X1   g119(.A(G113gat), .B(G141gat), .Z(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT91), .B(G197gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT11), .B(G169gat), .Z(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n314), .A3(new_n320), .A4(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n309), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n319), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n306), .A2(new_n313), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT109), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n256), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  XOR2_X1   g139(.A(G57gat), .B(G64gat), .Z(new_n341));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n342));
  INV_X1    g141(.A(G71gat), .ZN(new_n343));
  INV_X1    g142(.A(G78gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G71gat), .B(G78gat), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n345), .A3(new_n341), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n254), .A2(new_n338), .A3(new_n255), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n340), .A2(new_n348), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n350), .A2(new_n348), .A3(KEYINPUT105), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT105), .B1(new_n350), .B2(new_n348), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n258), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OR4_X1    g156(.A1(new_n356), .A2(new_n353), .A3(new_n258), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n337), .B1(new_n359), .B2(KEYINPUT110), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT110), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n352), .A2(new_n355), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n337), .ZN(new_n365));
  XNOR2_X1  g164(.A(G120gat), .B(G148gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G176gat), .B(G204gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n359), .A2(new_n336), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n335), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n300), .A2(KEYINPUT21), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n353), .B2(new_n354), .ZN(new_n377));
  XOR2_X1   g176(.A(G127gat), .B(G155gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G231gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(G183gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G211gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n379), .B(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n300), .A2(KEYINPUT21), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n384), .B(new_n387), .Z(new_n388));
  NAND3_X1  g187(.A1(new_n288), .A2(new_n375), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G190gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G169gat), .ZN(new_n394));
  INV_X1    g193(.A(G176gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT26), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT26), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n390), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT67), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n390), .C1(new_n400), .C2(new_n401), .ZN(new_n407));
  AOI211_X1 g206(.A(new_n391), .B(new_n399), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  AND3_X1   g208(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT23), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(G169gat), .B2(G176gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n416), .A3(new_n392), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n409), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT25), .ZN(new_n420));
  AND3_X1   g219(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n413), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n418), .A2(new_n419), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT65), .B(new_n409), .C1(new_n413), .C2(new_n417), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n408), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT77), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n419), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n396), .A2(new_n398), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n391), .B1(new_n434), .B2(new_n392), .ZN(new_n435));
  INV_X1    g234(.A(new_n407), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT27), .B(G183gat), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n404), .B1(new_n437), .B2(new_n390), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT77), .ZN(new_n441));
  INV_X1    g240(.A(new_n429), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(KEYINPUT68), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n406), .A2(new_n407), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n435), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n449), .B2(new_n433), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n430), .B(new_n443), .C1(new_n442), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT75), .B(G211gat), .ZN(new_n453));
  INV_X1    g252(.A(G218gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G211gat), .B(G218gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n445), .A2(new_n448), .B1(new_n426), .B2(new_n427), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n442), .A2(KEYINPUT29), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n466), .A2(new_n442), .B1(new_n440), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT78), .B1(new_n468), .B2(new_n464), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n467), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n433), .A3(new_n442), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n463), .ZN(new_n474));
  XNOR2_X1  g273(.A(G8gat), .B(G36gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n465), .A2(new_n469), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n473), .B1(new_n472), .B2(new_n463), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT78), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(KEYINPUT30), .A3(new_n465), .A4(new_n478), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  AND4_X1   g285(.A1(KEYINPUT79), .A2(new_n465), .A3(new_n469), .A4(new_n474), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT79), .B1(new_n484), .B2(new_n465), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n477), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(new_n248), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT0), .B(G57gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(G148gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G141gat), .ZN(new_n496));
  INV_X1    g295(.A(G141gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G148gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G141gat), .B(G148gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT2), .ZN(new_n503));
  INV_X1    g302(.A(G155gat), .ZN(new_n504));
  INV_X1    g303(.A(G162gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G155gat), .A2(G162gat), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n502), .A2(KEYINPUT81), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n503), .A2(KEYINPUT80), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n503), .A2(KEYINPUT80), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G155gat), .B(G162gat), .Z(new_n512));
  AOI22_X1  g311(.A1(new_n501), .A2(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G113gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(G120gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(G120gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(KEYINPUT71), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(KEYINPUT71), .B2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(G127gat), .ZN(new_n519));
  INV_X1    g318(.A(G134gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G127gat), .A2(G134gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT1), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT1), .ZN(new_n525));
  INV_X1    g324(.A(G120gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G113gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n515), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  NOR2_X1   g328(.A1(G127gat), .A2(G134gat), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT69), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n521), .B2(new_n522), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n528), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT69), .B1(new_n529), .B2(new_n530), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n532), .A3(new_n522), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n539), .B2(new_n528), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n513), .B(new_n524), .C1(new_n535), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n536), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n513), .A4(new_n524), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G225gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n502), .A2(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n506), .A2(new_n507), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n501), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT3), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n512), .B1(new_n502), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n552), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n524), .B1(new_n535), .B2(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n548), .A2(KEYINPUT5), .A3(new_n549), .A4(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n549), .ZN(new_n562));
  AOI221_X4 g361(.A(new_n562), .B1(new_n558), .B2(new_n559), .C1(new_n542), .C2(new_n547), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT5), .ZN(new_n564));
  INV_X1    g363(.A(new_n513), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n541), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n494), .B(new_n561), .C1(new_n563), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT6), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n543), .A2(new_n544), .B1(new_n518), .B2(new_n523), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n513), .ZN(new_n573));
  INV_X1    g372(.A(new_n541), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n562), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT5), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n549), .A3(new_n560), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n494), .B1(new_n578), .B2(new_n561), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n569), .B(new_n571), .C1(new_n579), .C2(KEYINPUT6), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n561), .B1(new_n563), .B2(new_n568), .ZN(new_n581));
  INV_X1    g380(.A(new_n494), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT6), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n569), .A2(new_n571), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT83), .B1(new_n490), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n465), .A2(new_n469), .A3(new_n474), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n484), .A2(KEYINPUT79), .A3(new_n465), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n478), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n481), .A2(new_n485), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n586), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT83), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n444), .B1(new_n460), .B2(new_n462), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n565), .B1(new_n599), .B2(KEYINPUT3), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n556), .A2(new_n444), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n464), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G228gat), .A2(G233gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n464), .B2(new_n601), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT29), .B1(new_n460), .B2(new_n462), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n565), .B1(new_n606), .B2(KEYINPUT3), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G22gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G78gat), .B(G106gat), .Z(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT85), .B(G50gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n603), .A2(new_n604), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n605), .A2(new_n607), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n609), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n608), .B2(new_n609), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n610), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n621), .A3(new_n615), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n608), .A2(new_n609), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT86), .B1(new_n608), .B2(new_n609), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n625), .B(new_n626), .C1(new_n615), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n448), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n447), .B1(new_n446), .B2(new_n435), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n433), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n559), .ZN(new_n633));
  NAND2_X1  g432(.A1(G227gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT64), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n449), .A2(new_n572), .A3(new_n433), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT34), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G15gat), .B(G43gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G71gat), .B(G99gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  AOI21_X1  g443(.A(new_n636), .B1(new_n633), .B2(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT32), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n449), .A2(new_n572), .A3(new_n433), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n572), .B1(new_n449), .B2(new_n433), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n635), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n653));
  INV_X1    g452(.A(new_n644), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n652), .B(KEYINPUT32), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n641), .B1(new_n649), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(KEYINPUT32), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n644), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n640), .A3(new_n655), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n657), .B1(KEYINPUT74), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT74), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n640), .B1(new_n655), .B2(new_n660), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT36), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT72), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n660), .A2(new_n667), .A3(new_n655), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n660), .B2(new_n655), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n641), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT73), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT73), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n672), .B(new_n641), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n671), .A2(KEYINPUT36), .A3(new_n661), .A4(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n598), .A2(new_n629), .B1(new_n666), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n588), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n477), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n451), .A2(new_n463), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT37), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n472), .B2(new_n464), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n465), .A2(new_n680), .A3(new_n469), .A4(new_n474), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n676), .A2(new_n478), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n586), .A2(KEYINPUT89), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT89), .B1(new_n586), .B2(new_n684), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT37), .B1(new_n487), .B2(new_n488), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n683), .A2(new_n477), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n677), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n548), .A2(new_n560), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n549), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT39), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n494), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n566), .A2(new_n549), .A3(new_n541), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(KEYINPUT88), .ZN(new_n696));
  OAI221_X1 g495(.A(new_n696), .B1(KEYINPUT88), .B2(new_n695), .C1(new_n691), .C2(new_n549), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n694), .A2(KEYINPUT40), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT40), .B1(new_n694), .B2(new_n697), .ZN(new_n699));
  INV_X1    g498(.A(new_n569), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n490), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n624), .A2(new_n628), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT90), .B1(new_n690), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n686), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n586), .A2(KEYINPUT89), .A3(new_n684), .ZN(new_n707));
  INV_X1    g506(.A(new_n689), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT90), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n629), .B1(new_n701), .B2(new_n490), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n675), .A2(new_n705), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n671), .A2(new_n703), .A3(new_n661), .A4(new_n673), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT35), .B1(new_n598), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n703), .B1(new_n662), .B2(new_n665), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT35), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n594), .A2(new_n595), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n389), .B1(new_n713), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n586), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g523(.A1(new_n722), .A2(new_n490), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n297), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT16), .B(G8gat), .Z(new_n727));
  AND2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT111), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(KEYINPUT42), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT42), .B2(new_n729), .ZN(G1325gat));
  INV_X1    g530(.A(new_n662), .ZN(new_n732));
  INV_X1    g531(.A(new_n665), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(G15gat), .B1(new_n722), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n666), .A2(new_n674), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT112), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(G15gat), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n722), .B2(new_n739), .ZN(G1326gat));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n629), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  AOI21_X1  g542(.A(new_n288), .B1(new_n713), .B2(new_n721), .ZN(new_n744));
  INV_X1    g543(.A(new_n388), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n375), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n586), .A3(new_n209), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n752), .B(new_n288), .C1(new_n713), .C2(new_n721), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n673), .A2(new_n661), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT72), .B1(new_n649), .B2(new_n656), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n660), .A2(new_n667), .A3(new_n655), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n672), .B1(new_n757), .B2(new_n641), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(new_n703), .A3(new_n587), .A4(new_n597), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT113), .B(new_n719), .C1(new_n760), .C2(KEYINPUT35), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n715), .B2(new_n720), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n713), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n283), .A2(new_n287), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n753), .B1(new_n766), .B2(new_n752), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n767), .B2(new_n747), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT44), .B1(new_n764), .B2(new_n765), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n770), .A2(new_n753), .A3(new_n771), .A4(new_n746), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n595), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n751), .B1(new_n774), .B2(new_n209), .ZN(G1328gat));
  NOR3_X1   g574(.A1(new_n748), .A2(G36gat), .A3(new_n594), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT46), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n594), .B1(new_n769), .B2(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n210), .ZN(G1329gat));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n747), .ZN(new_n780));
  OAI21_X1  g579(.A(G43gat), .B1(new_n780), .B2(new_n736), .ZN(new_n781));
  INV_X1    g580(.A(new_n734), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(G43gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n749), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  INV_X1    g584(.A(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n748), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n781), .A2(KEYINPUT47), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n788), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n738), .B1(new_n768), .B2(new_n772), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(G43gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g592(.A(G50gat), .B1(new_n780), .B2(new_n703), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n748), .A2(G50gat), .A3(new_n703), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(KEYINPUT48), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n629), .B1(new_n768), .B2(new_n772), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n798), .B2(G50gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g599(.A(new_n374), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n765), .A2(new_n334), .A3(new_n801), .A4(new_n745), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n764), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n586), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n594), .ZN(new_n807));
  NOR2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  AND2_X1   g607(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n807), .B2(new_n808), .ZN(G1333gat));
  OAI21_X1  g610(.A(new_n343), .B1(new_n803), .B2(new_n782), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n738), .A2(G71gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n803), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g614(.A1(new_n803), .A2(new_n703), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(new_n344), .ZN(G1335gat));
  NOR2_X1   g616(.A1(new_n388), .A2(new_n334), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n764), .A2(new_n765), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n764), .A2(new_n821), .A3(new_n765), .A4(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n374), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(new_n595), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n818), .A2(new_n374), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n770), .A2(new_n753), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n595), .A2(new_n248), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n824), .A2(new_n248), .B1(new_n826), .B2(new_n827), .ZN(G1336gat));
  AND2_X1   g627(.A1(new_n826), .A2(new_n490), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n490), .A2(new_n249), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n829), .A2(new_n249), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833));
  OAI221_X1 g632(.A(new_n833), .B1(new_n823), .B2(new_n830), .C1(new_n829), .C2(new_n249), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1337gat));
  NOR2_X1   g634(.A1(new_n782), .A2(G99gat), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n374), .A3(new_n822), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n721), .A2(KEYINPUT113), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n715), .A2(new_n762), .A3(new_n720), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n690), .A2(new_n704), .A3(KEYINPUT90), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n675), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n752), .B1(new_n843), .B2(new_n288), .ZN(new_n844));
  INV_X1    g643(.A(new_n753), .ZN(new_n845));
  INV_X1    g644(.A(new_n825), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n844), .A2(new_n738), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  OAI21_X1  g647(.A(G99gat), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT116), .B1(new_n826), .B2(new_n738), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n837), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1338gat));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n820), .A2(new_n629), .A3(new_n374), .A4(new_n822), .ZN(new_n858));
  INV_X1    g657(.A(G106gat), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n703), .A2(new_n859), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n826), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n856), .B(new_n857), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n858), .A2(new_n859), .B1(new_n826), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n864), .B2(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1339gat));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n307), .A2(new_n309), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n325), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n327), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n359), .A2(new_n873), .A3(new_n336), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n368), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n363), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT54), .B1(new_n359), .B2(new_n336), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n876), .B(KEYINPUT55), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n360), .B2(new_n362), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n875), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n879), .A2(new_n370), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n872), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n327), .A2(new_n871), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n884), .A2(new_n287), .A3(new_n283), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n334), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n327), .A2(new_n374), .A3(new_n871), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n288), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n388), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n288), .A2(new_n335), .A3(new_n801), .A4(new_n388), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n867), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n883), .A3(new_n872), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n288), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n888), .A2(new_n889), .B1(new_n283), .B2(new_n287), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n745), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT120), .A3(new_n893), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n716), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n490), .A2(new_n595), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G113gat), .B1(new_n904), .B2(new_n335), .ZN(new_n905));
  INV_X1    g704(.A(new_n714), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n334), .A2(new_n514), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1340gat));
  OAI21_X1  g708(.A(G120gat), .B1(new_n904), .B2(new_n801), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n374), .A2(new_n526), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n907), .B2(new_n911), .ZN(G1341gat));
  OAI21_X1  g711(.A(G127gat), .B1(new_n904), .B2(new_n745), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n388), .A2(new_n519), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT121), .ZN(G1342gat));
  NAND2_X1  g715(.A1(new_n765), .A2(new_n520), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n907), .A2(KEYINPUT56), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G134gat), .B1(new_n904), .B2(new_n288), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT56), .B1(new_n907), .B2(new_n917), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G1343gat));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n900), .A3(new_n629), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n736), .A2(new_n903), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n629), .B1(new_n892), .B2(new_n894), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n923), .A2(new_n334), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G141gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n922), .A2(new_n738), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n929), .A2(new_n497), .A3(new_n334), .A4(new_n903), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1344gat));
  NAND3_X1  g734(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n801), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G148gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n703), .A2(KEYINPUT57), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n897), .A2(new_n898), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT122), .B1(new_n887), .B2(new_n891), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n388), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n946), .B2(new_n894), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n374), .A3(new_n924), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n938), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n903), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n374), .A2(new_n495), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n940), .A2(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1345gat));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n504), .A3(new_n745), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n929), .A2(new_n388), .A3(new_n903), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n504), .ZN(G1346gat));
  NAND4_X1  g755(.A1(new_n923), .A2(new_n765), .A3(new_n924), .A4(new_n926), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT123), .ZN(new_n958));
  OAI21_X1  g757(.A(G162gat), .B1(new_n957), .B2(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n765), .A2(new_n505), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n958), .A2(new_n959), .B1(new_n951), .B2(new_n960), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n594), .A2(new_n586), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n895), .A2(new_n900), .A3(new_n902), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n335), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n901), .A2(new_n906), .A3(new_n962), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n334), .A2(new_n394), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1348gat));
  NOR3_X1   g766(.A1(new_n963), .A2(new_n395), .A3(new_n801), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n965), .A2(new_n801), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n395), .ZN(G1349gat));
  OR3_X1    g769(.A1(new_n963), .A2(KEYINPUT124), .A3(new_n745), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT124), .B1(new_n963), .B2(new_n745), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(G183gat), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n388), .A2(new_n437), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT60), .ZN(G1350gat));
  OR3_X1    g776(.A1(new_n965), .A2(G190gat), .A3(new_n288), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n963), .A2(new_n288), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(G190gat), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n979), .B(G190gat), .C1(new_n963), .C2(new_n288), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n978), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n978), .B(KEYINPUT125), .C1(new_n981), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1351gat));
  INV_X1    g787(.A(new_n962), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n738), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n948), .A2(new_n334), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G197gat), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n922), .A2(new_n738), .A3(new_n989), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n335), .A2(G197gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1352gat));
  INV_X1    g795(.A(G204gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n374), .A2(new_n997), .ZN(new_n998));
  OR3_X1    g797(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT62), .B1(new_n994), .B2(new_n998), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n948), .A2(new_n374), .A3(new_n990), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n999), .B(new_n1000), .C1(new_n1001), .C2(new_n997), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n993), .A2(new_n453), .A3(new_n388), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n941), .A2(new_n388), .A3(new_n947), .A4(new_n990), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G211gat), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  OAI21_X1  g811(.A(new_n454), .B1(new_n994), .B2(new_n288), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n288), .A2(new_n454), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n948), .A2(new_n990), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1013), .A2(new_n1015), .A3(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(G1355gat));
endmodule


