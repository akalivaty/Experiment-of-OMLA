//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT94), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(KEYINPUT16), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(G8gat), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT95), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n203), .A2(KEYINPUT95), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n212), .C1(new_n208), .C2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220));
  OR3_X1    g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n219), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n218), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n225), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT17), .B1(new_n225), .B2(KEYINPUT93), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n215), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n225), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(KEYINPUT13), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n231), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n230), .A2(new_n225), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n240), .A2(KEYINPUT96), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT96), .B1(new_n240), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n239), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G113gat), .B(G141gat), .Z(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n244), .A2(KEYINPUT97), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT97), .B1(new_n244), .B2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n241), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n256), .B2(new_n238), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G22gat), .B(G50gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G141gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G148gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT78), .B(G148gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT2), .ZN(new_n267));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT80), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(new_n271), .A3(new_n267), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G148gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G141gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n268), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284));
  INV_X1    g083(.A(G211gat), .ZN(new_n285));
  INV_X1    g084(.A(G218gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n282), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n282), .B(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n283), .A2(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT29), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n281), .B1(new_n296), .B2(KEYINPUT3), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT88), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n295), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(KEYINPUT88), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G228gat), .A3(G233gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n306), .B(KEYINPUT31), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n270), .A2(new_n272), .B1(new_n279), .B2(new_n278), .ZN(new_n310));
  INV_X1    g109(.A(new_n292), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n290), .B1(new_n282), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT3), .B1(new_n312), .B2(new_n300), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n302), .B(new_n309), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n308), .B1(new_n305), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n261), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n260), .A3(new_n315), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT81), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G113gat), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT69), .B(G120gat), .Z(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(G113gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n328), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT69), .B(G120gat), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(new_n336), .B2(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n324), .A2(KEYINPUT67), .A3(new_n325), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n335), .A2(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n328), .B2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n339), .A2(new_n342), .A3(KEYINPUT68), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n322), .B1(new_n281), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n332), .A2(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n310), .A2(new_n351), .A3(KEYINPUT81), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n281), .A2(new_n349), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT83), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n350), .A2(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n299), .A2(new_n349), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n281), .A2(new_n349), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT4), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n363), .A2(new_n355), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(new_n369), .A3(new_n358), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n360), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n358), .A2(new_n356), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n310), .A2(new_n351), .A3(new_n362), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT84), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n350), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n366), .A2(KEYINPUT84), .A3(new_n362), .ZN(new_n380));
  AND4_X1   g179(.A1(new_n373), .A2(new_n376), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n372), .B(new_n365), .C1(new_n377), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT0), .B(G57gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G85gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n382), .A3(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT86), .B1(new_n390), .B2(new_n391), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397));
  INV_X1    g196(.A(G64gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(G92gat), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G226gat), .ZN(new_n402));
  INV_X1    g201(.A(G233gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT24), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(G183gat), .B2(G190gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT23), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n409), .A2(KEYINPUT23), .ZN(new_n411));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT66), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n408), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(KEYINPUT66), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT25), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n410), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n417), .B2(KEYINPUT65), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(KEYINPUT65), .B2(new_n417), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT25), .ZN(new_n420));
  NOR2_X1   g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT64), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n407), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n419), .A2(new_n420), .A3(new_n411), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT27), .B(G183gat), .ZN(new_n425));
  INV_X1    g224(.A(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT28), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT26), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n412), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n406), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n424), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n416), .A2(new_n424), .A3(KEYINPUT74), .A4(new_n434), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n405), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n404), .A2(KEYINPUT29), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n439), .A2(new_n441), .A3(new_n294), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n435), .A2(new_n405), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n295), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NOR4_X1   g246(.A1(new_n439), .A2(KEYINPUT75), .A3(new_n441), .A4(new_n294), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n401), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n445), .A2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(new_n442), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n448), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n400), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n449), .B2(new_n451), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n453), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT87), .B1(new_n396), .B2(new_n460), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n321), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n365), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n375), .A2(new_n376), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT85), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n375), .A2(new_n373), .A3(new_n376), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OR3_X1    g267(.A1(new_n468), .A2(KEYINPUT39), .A3(new_n355), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n361), .A2(new_n355), .A3(new_n353), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT39), .B(new_n470), .C1(new_n468), .C2(new_n355), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n387), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n456), .A2(new_n400), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT76), .B1(new_n475), .B2(KEYINPUT30), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(KEYINPUT30), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n457), .A4(new_n452), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n383), .B2(new_n388), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n383), .A2(new_n479), .A3(new_n388), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n472), .A2(new_n473), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n474), .A2(new_n478), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n318), .A2(new_n320), .ZN(new_n486));
  INV_X1    g285(.A(new_n482), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n391), .B(new_n390), .C1(new_n487), .C2(new_n480), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n456), .A2(KEYINPUT37), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n401), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n439), .A2(new_n441), .A3(new_n295), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n294), .B1(new_n443), .B2(new_n444), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n389), .A3(new_n449), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n456), .A2(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n491), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n485), .B(new_n486), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n435), .B(new_n351), .ZN(new_n504));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n506), .B2(KEYINPUT33), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n504), .A2(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n507), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT32), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n511), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT36), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n463), .A2(new_n500), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n396), .A2(new_n460), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n460), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n486), .A2(new_n515), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n390), .A2(new_n391), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n481), .B2(new_n482), .ZN(new_n526));
  INV_X1    g325(.A(new_n389), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n460), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n528), .B2(KEYINPUT90), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n478), .B1(new_n488), .B2(new_n389), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT35), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n524), .A2(KEYINPUT35), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT91), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n463), .A2(new_n500), .A3(new_n516), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n259), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n398), .A2(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n546), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n215), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G183gat), .ZN(new_n558));
  INV_X1    g357(.A(G183gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n215), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n558), .B2(new_n560), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n285), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n563), .B2(new_n564), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n567), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  AND2_X1   g380(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT8), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n579), .A2(new_n580), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT8), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(G99gat), .B2(G106gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT100), .B(G92gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(new_n581), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n580), .B1(new_n593), .B2(new_n579), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n596));
  INV_X1    g395(.A(new_n580), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n596), .A2(KEYINPUT101), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n226), .B2(new_n227), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n588), .A3(new_n587), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n589), .A2(new_n594), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n225), .ZN(new_n605));
  NAND3_X1  g404(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT102), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT98), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n607), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n607), .B2(new_n610), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n616), .B2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT108), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G120gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n274), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n555), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n555), .A2(new_n601), .A3(new_n587), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n555), .A2(new_n601), .A3(KEYINPUT104), .A4(new_n587), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n599), .A2(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n547), .A2(new_n554), .A3(KEYINPUT10), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n595), .B2(new_n598), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT106), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n604), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n602), .A2(new_n603), .A3(new_n629), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT107), .B1(new_n645), .B2(new_n628), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647));
  INV_X1    g446(.A(new_n628), .ZN(new_n648));
  AOI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n640), .C2(new_n644), .ZN(new_n649));
  OAI221_X1 g448(.A(new_n627), .B1(new_n628), .B2(new_n634), .C1(new_n646), .C2(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n634), .A2(new_n643), .B1(new_n637), .B2(new_n639), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n648), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n634), .A2(new_n628), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n626), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n574), .A2(new_n622), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n541), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n396), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n207), .ZN(G1324gat));
  NAND3_X1  g458(.A1(new_n541), .A2(new_n478), .A3(new_n656), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n660), .A2(new_n666), .A3(G8gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n660), .B2(G8gat), .ZN(new_n668));
  OAI22_X1  g467(.A1(new_n664), .A2(new_n665), .B1(new_n667), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n657), .A2(new_n670), .A3(new_n516), .ZN(new_n671));
  INV_X1    g470(.A(new_n515), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n657), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(KEYINPUT110), .B(new_n670), .C1(new_n657), .C2(new_n672), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n657), .A2(new_n486), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n534), .A2(new_n540), .ZN(new_n681));
  INV_X1    g480(.A(new_n622), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n622), .B1(new_n517), .B2(new_n533), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n681), .A2(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n574), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n655), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n258), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n396), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n687), .A2(new_n682), .A3(new_n655), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n541), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n396), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR4_X1   g496(.A1(new_n694), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n396), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n690), .B1(new_n697), .B2(new_n698), .ZN(G1328gat));
  OAI21_X1  g498(.A(G36gat), .B1(new_n689), .B2(new_n460), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n460), .A2(G36gat), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT46), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n694), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(G1329gat));
  INV_X1    g503(.A(G43gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n516), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n686), .A2(new_n258), .A3(new_n688), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n541), .A2(new_n515), .A3(new_n692), .A4(new_n693), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1330gat));
  INV_X1    g513(.A(G50gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n486), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n686), .A2(new_n258), .A3(new_n688), .A4(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n541), .A2(new_n321), .A3(new_n692), .A4(new_n693), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n715), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT48), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT48), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1331gat));
  INV_X1    g521(.A(new_n655), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n537), .B2(new_n539), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n258), .A2(new_n574), .A3(new_n622), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n396), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n548), .ZN(G1332gat));
  AOI211_X1 g527(.A(new_n460), .B(new_n726), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  OR3_X1    g530(.A1(new_n726), .A2(G71gat), .A3(new_n672), .ZN(new_n732));
  OAI21_X1  g531(.A(G71gat), .B1(new_n726), .B2(new_n516), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n726), .A2(new_n486), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g537(.A1(new_n258), .A2(new_n687), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n723), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n686), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(new_n581), .A3(new_n396), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n685), .B2(new_n740), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n537), .A2(new_n539), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(KEYINPUT51), .A3(new_n622), .A4(new_n739), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n746), .ZN(new_n750));
  INV_X1    g549(.A(new_n396), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .A4(new_n655), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n743), .B1(new_n581), .B2(new_n752), .ZN(G1336gat));
  NAND2_X1  g552(.A1(new_n681), .A2(new_n684), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n747), .B2(new_n622), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n754), .A2(new_n756), .A3(new_n478), .A4(new_n741), .ZN(new_n757));
  INV_X1    g556(.A(new_n592), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n460), .A2(G92gat), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n655), .A2(new_n749), .A3(new_n750), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n723), .B1(new_n745), .B2(new_n748), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n757), .A2(new_n758), .B1(new_n764), .B2(new_n762), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n761), .A2(new_n763), .B1(new_n765), .B2(new_n760), .ZN(G1337gat));
  XOR2_X1   g565(.A(KEYINPUT113), .B(G99gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n742), .B2(new_n516), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n672), .A2(new_n767), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n750), .A3(new_n655), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n756), .A3(new_n321), .A4(new_n741), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n486), .A2(G106gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n749), .A2(new_n750), .A3(new_n655), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n772), .A2(G106gat), .B1(new_n764), .B2(new_n774), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n651), .B2(new_n648), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n646), .B2(new_n649), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT115), .B(new_n783), .C1(new_n646), .C2(new_n649), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n652), .A2(new_n782), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n626), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n781), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(KEYINPUT55), .B(new_n790), .C1(new_n786), .C2(new_n787), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n650), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n235), .A2(new_n236), .A3(new_n234), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n228), .A2(new_n231), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n229), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n249), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n254), .A2(new_n622), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT116), .B(new_n650), .C1(new_n792), .C2(new_n793), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n796), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n796), .A2(new_n801), .A3(KEYINPUT117), .A4(new_n802), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n796), .A2(new_n258), .A3(new_n802), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n254), .A2(new_n655), .A3(new_n800), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n622), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n574), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n259), .A2(new_n656), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n522), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n751), .A2(new_n460), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n259), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(new_n335), .ZN(G1340gat));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n723), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n329), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n327), .B2(new_n819), .ZN(G1341gat));
  NOR2_X1   g620(.A1(new_n816), .A2(new_n574), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(G127gat), .Z(G1342gat));
  NAND3_X1  g622(.A1(new_n813), .A2(new_n622), .A3(new_n815), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n824), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(G134gat), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT56), .B1(new_n824), .B2(G134gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(G1343gat));
  AOI21_X1  g627(.A(new_n486), .B1(new_n811), .B2(new_n812), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT119), .A3(new_n751), .A4(new_n516), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n805), .A2(new_n806), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n808), .A2(new_n809), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n682), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n687), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n812), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n321), .B(new_n516), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(new_n396), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n478), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n259), .A2(G141gat), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n829), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n815), .A2(new_n516), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT118), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n809), .B1(new_n259), .B2(new_n794), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n682), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n687), .B1(new_n832), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n321), .B1(new_n848), .B2(new_n836), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT57), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n843), .A2(new_n258), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G141gat), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n516), .A2(new_n829), .A3(new_n815), .A4(new_n840), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n851), .B2(G141gat), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n841), .A2(new_n854), .B1(new_n853), .B2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n274), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n812), .B(KEYINPUT120), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n254), .A2(new_n622), .A3(new_n800), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n794), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n846), .B2(new_n682), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n860), .B1(new_n687), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n321), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n842), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n829), .A2(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n655), .A3(new_n845), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n843), .A2(new_n845), .A3(new_n850), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(KEYINPUT59), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n859), .A2(new_n872), .B1(new_n874), .B2(new_n655), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n858), .B1(new_n839), .B2(new_n655), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n264), .B2(new_n876), .ZN(G1345gat));
  XNOR2_X1  g676(.A(KEYINPUT79), .B(G155gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n839), .B2(new_n687), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n873), .A2(new_n574), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(G1346gat));
  OAI21_X1  g680(.A(G162gat), .B1(new_n873), .B2(new_n682), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n478), .B(new_n682), .C1(new_n830), .C2(new_n838), .ZN(new_n883));
  INV_X1    g682(.A(G162gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT122), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n830), .A2(new_n838), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n884), .A3(new_n460), .A4(new_n622), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n882), .B1(new_n885), .B2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n751), .A2(new_n460), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n813), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n259), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT124), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n813), .A2(KEYINPUT123), .A3(new_n891), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G169gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n258), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n900), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n898), .B2(new_n655), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n892), .A2(new_n723), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(G176gat), .B2(new_n903), .ZN(G1349gat));
  NOR2_X1   g703(.A1(new_n892), .A2(new_n574), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n425), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n905), .B2(new_n559), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n906), .B(new_n909), .C1(new_n559), .C2(new_n905), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n892), .B2(new_n682), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT61), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n426), .A3(new_n622), .A4(new_n897), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n891), .A2(new_n516), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n871), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n259), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n829), .A2(new_n920), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n923), .A2(G197gat), .A3(new_n259), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1352gat));
  NOR3_X1   g724(.A1(new_n923), .A2(G204gat), .A3(new_n723), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n927), .B2(KEYINPUT62), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n921), .B2(new_n723), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(new_n923), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n285), .A3(new_n687), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n871), .A2(new_n687), .A3(new_n920), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  NAND2_X1  g739(.A1(new_n622), .A2(G218gat), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT127), .Z(new_n942));
  NOR2_X1   g741(.A1(new_n921), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G218gat), .B1(new_n935), .B2(new_n622), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


