//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT67), .B(G244), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n212), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n213), .C2(new_n214), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT64), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n228), .B1(new_n202), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n230), .B1(new_n229), .B2(new_n202), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n210), .B(new_n224), .C1(new_n227), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT69), .B(G50), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  AND3_X1   g0050(.A1(new_n250), .A2(KEYINPUT70), .A3(new_n225), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT70), .B1(new_n250), .B2(new_n225), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT72), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n254), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G50), .B2(new_n267), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n276), .B1(new_n216), .B2(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G200), .B2(new_n291), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n272), .A2(new_n273), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(new_n291), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n270), .B1(new_n297), .B2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n291), .A2(G179), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n274), .A2(G226), .A3(new_n275), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n283), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  INV_X1    g0108(.A(new_n287), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n285), .A2(KEYINPUT74), .A3(new_n286), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n311), .B1(new_n289), .B2(G238), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n307), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n308), .B1(new_n312), .B2(new_n307), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT14), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(G169), .C1(new_n313), .C2(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(G179), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n260), .A2(G50), .ZN(new_n322));
  INV_X1    g0122(.A(new_n258), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n322), .B1(new_n226), .B2(G68), .C1(new_n216), .C2(new_n323), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n253), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n250), .A2(new_n225), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G68), .A3(new_n264), .ZN(new_n328));
  INV_X1    g0128(.A(new_n267), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT12), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT12), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n267), .B2(G68), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n326), .A2(new_n328), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n325), .B1(new_n324), .B2(new_n253), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n321), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n315), .A2(G190), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n256), .A2(new_n264), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n343), .A2(new_n253), .B1(new_n267), .B2(new_n256), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n330), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n201), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n260), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(G33), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(G33), .ZN(new_n356));
  AOI21_X1  g0156(.A(G20), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT77), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT76), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n363), .A2(new_n358), .A3(new_n226), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n226), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n330), .B1(new_n366), .B2(KEYINPUT7), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n357), .A2(new_n358), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT77), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n350), .C1(new_n365), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n250), .A2(new_n225), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n358), .B1(new_n274), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n354), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n349), .B1(new_n376), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n371), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n344), .B1(new_n370), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n278), .A2(new_n275), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n275), .A2(G226), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n355), .A2(new_n356), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n282), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n309), .B1(new_n288), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n382), .A2(new_n381), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n384), .B1(new_n363), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n283), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT79), .B(G190), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n388), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n380), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT17), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n380), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n316), .B1(new_n385), .B2(new_n387), .ZN(new_n404));
  INV_X1    g0204(.A(G179), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n392), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n404), .B2(new_n406), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n403), .B1(new_n380), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n404), .A2(new_n406), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n408), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n360), .B1(new_n359), .B2(new_n364), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n368), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n349), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n378), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n415), .B(KEYINPUT18), .C1(new_n419), .C2(new_n344), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n402), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n309), .B1(new_n288), .B2(new_n217), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  INV_X1    g0226(.A(G238), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n425), .B1(new_n426), .B2(new_n274), .C1(new_n277), .C2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(new_n283), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n255), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n323), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(new_n371), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n327), .A2(G77), .A3(new_n264), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G77), .B2(new_n267), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n423), .B1(new_n429), .B2(G169), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n429), .A2(new_n405), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n433), .B2(new_n371), .ZN(new_n440));
  INV_X1    g0240(.A(new_n429), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(new_n316), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n423), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n429), .A2(G190), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n440), .C1(new_n446), .C2(new_n429), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR4_X1   g0248(.A1(new_n302), .A2(new_n342), .A3(new_n422), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n263), .B(G45), .C1(new_n452), .C2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT83), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n450), .A2(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(KEYINPUT83), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n283), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(KEYINPUT91), .A3(G264), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT91), .B1(new_n460), .B2(G264), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n263), .A2(G45), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n451), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n286), .B1(new_n280), .B2(new_n281), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n466), .A2(new_n459), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n455), .A2(new_n471), .A3(new_n459), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n221), .A2(G1698), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G250), .B2(G1698), .ZN(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n363), .A2(new_n475), .B1(new_n257), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n446), .B1(new_n463), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n460), .A2(G264), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n473), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n292), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n226), .A2(G87), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n374), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT23), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n226), .B2(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n426), .A2(KEYINPUT23), .A3(G20), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT88), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(G87), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n485), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n355), .A2(new_n226), .A3(new_n356), .A4(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n499), .A2(new_n496), .A3(new_n487), .A4(new_n493), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n487), .A3(new_n493), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT89), .B1(new_n505), .B2(new_n371), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(KEYINPUT89), .A3(new_n371), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n329), .A2(new_n426), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT90), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT25), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT81), .B1(new_n257), .B2(G1), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n263), .A3(G33), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n267), .B(new_n517), .C1(new_n251), .C2(new_n252), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n426), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n512), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n484), .A2(new_n507), .A3(new_n508), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n470), .A2(new_n472), .B1(new_n460), .B2(G257), .ZN(new_n523));
  AND2_X1   g0323(.A1(KEYINPUT4), .A2(G244), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n354), .A2(new_n373), .A3(new_n524), .A4(new_n275), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n274), .A2(KEYINPUT82), .A3(new_n275), .A4(new_n524), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n257), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n354), .B2(new_n353), .ZN(new_n533));
  INV_X1    g0333(.A(G244), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT4), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n283), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n523), .A2(new_n537), .A3(G190), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n267), .A2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n518), .B2(new_n220), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT7), .B1(new_n374), .B2(new_n226), .ZN(new_n542));
  AOI211_X1 g0342(.A(new_n358), .B(G20), .C1(new_n354), .C2(new_n373), .ZN(new_n543));
  OAI21_X1  g0343(.A(G107), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g0344(.A(KEYINPUT80), .B(G107), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n220), .A2(KEYINPUT6), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n220), .A2(new_n426), .A3(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n548), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(G20), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n260), .A2(G77), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n544), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n541), .B1(new_n554), .B2(new_n371), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n538), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n446), .B1(new_n523), .B2(new_n537), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n522), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n557), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n559), .A2(KEYINPUT85), .A3(new_n555), .A4(new_n538), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G238), .A2(G1698), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n534), .B2(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n355), .A2(new_n563), .A3(new_n356), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n282), .B1(new_n564), .B2(new_n488), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n465), .A2(G250), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n282), .B1(new_n457), .B2(G274), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n405), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n226), .B1(new_n305), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n497), .A2(new_n220), .A3(new_n426), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n573), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n355), .A2(new_n226), .A3(new_n356), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n330), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n371), .ZN(new_n578));
  INV_X1    g0378(.A(new_n518), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n431), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n432), .A2(new_n329), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n316), .B1(new_n565), .B2(new_n568), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n564), .A2(new_n488), .ZN(new_n585));
  OAI211_X1 g0385(.A(G190), .B(new_n567), .C1(new_n585), .C2(new_n282), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n577), .A2(new_n371), .B1(new_n329), .B2(new_n432), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n565), .B2(new_n568), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(G87), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n523), .A2(new_n537), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n316), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n523), .A2(new_n537), .A3(new_n405), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n554), .A2(new_n371), .ZN(new_n596));
  INV_X1    g0396(.A(new_n541), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n521), .A2(new_n561), .A3(new_n592), .A4(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n517), .A2(new_n327), .A3(G116), .A4(new_n267), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT86), .ZN(new_n602));
  INV_X1    g0402(.A(G116), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n329), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n327), .A4(new_n517), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n530), .B(new_n226), .C1(G33), .C2(new_n220), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(G20), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n371), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n267), .A2(G116), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n607), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n221), .A2(new_n275), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(G264), .B2(new_n275), .ZN(new_n617));
  INV_X1    g0417(.A(G303), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n363), .A2(new_n617), .B1(new_n618), .B2(new_n274), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n283), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n460), .A2(G270), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n473), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n615), .B1(new_n622), .B2(G200), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n621), .A2(new_n620), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n394), .A3(new_n473), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n615), .A3(G169), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n622), .A2(new_n615), .A3(KEYINPUT21), .A4(G169), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n624), .A2(new_n615), .A3(G179), .A4(new_n473), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n626), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n629), .A4(new_n626), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n507), .A2(new_n508), .A3(new_n520), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT91), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n481), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n460), .A2(KEYINPUT91), .A3(G264), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n473), .A3(new_n478), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n642), .A2(new_n405), .B1(new_n316), .B2(new_n482), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n633), .A2(new_n636), .B1(new_n637), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n449), .A2(new_n600), .A3(new_n644), .ZN(G372));
  AND3_X1   g0445(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n558), .B2(new_n560), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n521), .A3(new_n592), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n508), .A2(new_n520), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n649), .B2(new_n506), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n584), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n594), .A2(new_n598), .A3(new_n655), .A4(new_n595), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n592), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n592), .A2(new_n646), .A3(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n449), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n337), .A2(new_n444), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n402), .A3(new_n341), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n421), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n300), .B1(new_n668), .B2(new_n296), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n263), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n637), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n521), .A3(new_n650), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n637), .A2(new_n643), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n633), .A2(new_n636), .B1(new_n615), .B2(new_n678), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n615), .A2(new_n678), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n651), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n678), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n637), .A2(new_n643), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n651), .A2(new_n678), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n682), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n208), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n573), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n232), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n703), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n599), .A2(new_n591), .A3(KEYINPUT26), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n710), .B(new_n584), .C1(new_n648), .C2(new_n652), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n657), .A2(new_n659), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT93), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n661), .A3(new_n660), .ZN(new_n717));
  INV_X1    g0517(.A(new_n584), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n650), .A2(new_n651), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n600), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n678), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n712), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n714), .B1(new_n722), .B2(KEYINPUT95), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n644), .A2(new_n600), .A3(new_n695), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n641), .A2(new_n478), .A3(new_n569), .ZN(new_n726));
  INV_X1    g0526(.A(new_n593), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n622), .A2(new_n405), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n727), .A4(new_n728), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n569), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n642), .A2(new_n593), .A3(new_n622), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n725), .B1(new_n735), .B2(new_n678), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(new_n725), .A3(new_n678), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n708), .B1(new_n742), .B2(G1), .ZN(G364));
  XNOR2_X1  g0543(.A(new_n691), .B(KEYINPUT96), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n263), .B1(new_n672), .B2(G45), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n703), .A2(KEYINPUT97), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT97), .ZN(new_n747));
  INV_X1    g0547(.A(new_n745), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n702), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n689), .B2(new_n690), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n225), .B1(G20), .B2(new_n316), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT98), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT98), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(G20), .A2(G179), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT99), .Z(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G200), .A3(new_n394), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n226), .B1(new_n763), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n762), .A2(G326), .B1(G294), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n760), .A2(new_n292), .A3(new_n446), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT102), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n446), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G20), .A3(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n226), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n763), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G303), .B1(new_n776), .B2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n771), .A2(new_n774), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n374), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n760), .A2(new_n446), .A3(new_n394), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G322), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n760), .A2(new_n292), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT101), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT33), .B(G317), .Z(new_n789));
  OAI211_X1 g0589(.A(new_n770), .B(new_n783), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n764), .A2(new_n220), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n775), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT100), .B(KEYINPUT32), .Z(new_n794));
  XNOR2_X1  g0594(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n768), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n791), .B(new_n795), .C1(G77), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n773), .A2(G87), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n374), .B1(new_n799), .B2(G107), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(new_n761), .C2(new_n228), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G58), .B2(new_n782), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n797), .B(new_n802), .C1(new_n330), .C2(new_n788), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n758), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n757), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n274), .A2(G355), .A3(new_n208), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n533), .A2(new_n701), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n706), .B2(G45), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n245), .A2(new_n456), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(G116), .B2(new_n208), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n750), .B(new_n804), .C1(new_n808), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n689), .A2(new_n807), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n753), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n757), .A2(new_n805), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n750), .B1(new_n819), .B2(new_n216), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n788), .A2(new_n778), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n768), .A2(new_n603), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n274), .B1(new_n773), .B2(G107), .ZN(new_n823));
  INV_X1    g0623(.A(new_n791), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n799), .A2(G87), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n776), .A2(G311), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n476), .A2(new_n781), .B1(new_n761), .B2(new_n618), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n821), .A2(new_n822), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n799), .A2(G68), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n228), .B2(new_n772), .C1(new_n831), .C2(new_n775), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n533), .B1(new_n345), .B2(new_n764), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G137), .A2(new_n762), .B1(new_n782), .B2(G143), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n792), .B2(new_n768), .C1(new_n788), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n832), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n829), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT103), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n447), .C1(new_n439), .C2(new_n443), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n678), .B1(new_n434), .B2(new_n436), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n444), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n820), .B1(new_n758), .B2(new_n840), .C1(new_n848), .C2(new_n806), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n721), .A2(new_n848), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n678), .B(new_n847), .C1(new_n717), .C2(new_n720), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n750), .B1(new_n853), .B2(new_n740), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(KEYINPUT104), .B1(new_n741), .B2(new_n852), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n849), .B1(new_n855), .B2(new_n856), .ZN(G384));
  NOR3_X1   g0657(.A1(new_n706), .A2(new_n216), .A3(new_n346), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n330), .A2(G50), .ZN(new_n859));
  OAI211_X1 g0659(.A(G1), .B(new_n671), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n550), .A2(new_n551), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n550), .A2(KEYINPUT35), .A3(new_n551), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(G116), .A4(new_n227), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  INV_X1    g0666(.A(new_n669), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n723), .B2(new_n449), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT107), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT106), .ZN(new_n870));
  INV_X1    g0670(.A(new_n676), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n421), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n337), .B(new_n341), .C1(new_n339), .C2(new_n695), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n321), .A2(new_n336), .A3(new_n678), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n444), .A2(new_n678), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n851), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n370), .A2(new_n379), .ZN(new_n879));
  INV_X1    g0679(.A(new_n344), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n879), .A2(new_n880), .B1(new_n414), .B2(new_n408), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n344), .B(new_n396), .C1(new_n370), .C2(new_n379), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n871), .B1(new_n419), .B2(new_n344), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT105), .B(new_n253), .C1(new_n418), .C2(KEYINPUT16), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n370), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n350), .B1(new_n365), .B2(new_n369), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT16), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT105), .B1(new_n891), .B2(new_n253), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n880), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n415), .A2(new_n871), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n882), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n886), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  INV_X1    g0697(.A(new_n370), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n254), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(KEYINPUT105), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n253), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n344), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n676), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n422), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n897), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n873), .B1(new_n878), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n337), .A2(new_n678), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n415), .B1(new_n419), .B2(new_n344), .ZN(new_n916));
  AND4_X1   g0716(.A1(new_n884), .A2(new_n916), .A3(new_n885), .A4(new_n398), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n399), .A2(new_n401), .B1(new_n412), .B2(new_n420), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n915), .A2(new_n917), .B1(new_n918), .B2(new_n885), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n912), .B1(new_n913), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n870), .B1(new_n910), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n398), .B1(new_n904), .B2(new_n894), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n917), .B1(new_n926), .B2(KEYINPUT37), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n918), .A2(new_n676), .A3(new_n904), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n920), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n922), .B1(new_n929), .B2(new_n914), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n914), .A2(new_n922), .A3(new_n921), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n911), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n876), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n695), .B(new_n848), .C1(new_n664), .C2(new_n653), .ZN(new_n934));
  INV_X1    g0734(.A(new_n877), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n929), .A2(new_n914), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n872), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n932), .A2(new_n938), .A3(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n869), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n847), .B1(new_n875), .B2(new_n874), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n739), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n914), .A2(new_n921), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n937), .A2(new_n739), .A3(new_n942), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n945), .A2(new_n946), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(G330), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n741), .A2(new_n449), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n449), .A2(new_n739), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n941), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n941), .A2(new_n952), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n953), .B1(new_n263), .B2(new_n672), .C1(new_n954), .C2(KEYINPUT108), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n860), .B(new_n866), .C1(new_n955), .C2(new_n956), .ZN(G367));
  AOI21_X1  g0757(.A(new_n374), .B1(new_n773), .B2(G58), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n799), .A2(G77), .ZN(new_n959));
  INV_X1    g0759(.A(G137), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n775), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G143), .B2(new_n762), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n228), .B2(new_n768), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT112), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n765), .A2(G68), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n781), .B2(new_n835), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n964), .B2(new_n966), .C1(new_n792), .C2(new_n788), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n788), .A2(new_n476), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n772), .B2(new_n603), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(new_n426), .C2(new_n764), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G283), .B2(new_n796), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n799), .A2(G97), .ZN(new_n975));
  INV_X1    g0775(.A(G317), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n363), .C1(new_n976), .C2(new_n775), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G303), .B2(new_n782), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(new_n767), .C2(new_n761), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n968), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT47), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n758), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n587), .A2(new_n589), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n678), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n592), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n584), .A2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n807), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n808), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n240), .A2(new_n701), .A3(new_n533), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n701), .C2(new_n431), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n751), .B1(new_n991), .B2(KEYINPUT111), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(KEYINPUT111), .B2(new_n991), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(new_n988), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n647), .B1(new_n555), .B2(new_n695), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n646), .A2(new_n678), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n698), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT44), .Z(new_n1001));
  OAI211_X1 g0801(.A(new_n696), .B(new_n998), .C1(new_n682), .C2(new_n697), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n693), .A2(KEYINPUT109), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT109), .B(new_n693), .C1(new_n1007), .C2(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n682), .A2(new_n683), .A3(new_n697), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n682), .A2(new_n697), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT110), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n682), .A2(new_n1014), .A3(new_n683), .A4(new_n697), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n692), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n744), .B2(new_n1016), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n741), .B(new_n723), .C1(new_n1010), .C2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n702), .B(KEYINPUT41), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n745), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1013), .A2(new_n996), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(KEYINPUT42), .B1(new_n646), .B2(new_n695), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n699), .A2(new_n996), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n986), .A2(new_n987), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1024), .A2(new_n1026), .B1(KEYINPUT43), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n694), .A2(new_n999), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n995), .B1(new_n1022), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n685), .A2(new_n807), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n810), .B1(new_n237), .B2(new_n456), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n274), .A2(new_n208), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n704), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n255), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n1042), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n1042), .B2(G50), .ZN(new_n1044));
  AOI21_X1  g0844(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1043), .A2(new_n704), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1041), .A2(new_n1046), .B1(new_n426), .B2(new_n701), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n751), .B1(new_n1047), .B2(new_n989), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n788), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n256), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n228), .A2(new_n781), .B1(new_n761), .B2(new_n792), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n773), .A2(G77), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n975), .C1(new_n835), .C2(new_n775), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n432), .A2(new_n764), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1053), .A3(new_n363), .A4(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1050), .B(new_n1055), .C1(new_n330), .C2(new_n768), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n799), .A2(G116), .B1(new_n776), .B2(G326), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n782), .B1(new_n762), .B2(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n618), .B2(new_n768), .C1(new_n788), .C2(new_n767), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT48), .Z(new_n1060));
  OAI22_X1  g0860(.A1(new_n772), .A2(new_n476), .B1(new_n764), .B2(new_n778), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n363), .B(new_n1057), .C1(new_n1062), .C2(KEYINPUT49), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n757), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1018), .A2(new_n748), .B1(new_n1038), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1018), .A2(new_n742), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n702), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1018), .A2(new_n742), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  OAI21_X1  g0871(.A(new_n702), .B1(new_n1009), .B2(new_n1068), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT116), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1001), .A2(new_n1004), .A3(new_n694), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n693), .B1(new_n1007), .B2(new_n1003), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1068), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1073), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT116), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n248), .A2(new_n810), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n808), .B1(new_n220), .B2(new_n208), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n788), .A2(new_n228), .B1(new_n1042), .B2(new_n768), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n835), .A2(new_n761), .B1(new_n781), .B2(new_n792), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT51), .Z(new_n1088));
  NAND2_X1  g0888(.A1(new_n776), .A2(G143), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n825), .B(new_n1089), .C1(new_n330), .C2(new_n772), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n533), .B1(new_n216), .B2(new_n764), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n274), .B1(new_n799), .B2(G107), .ZN(new_n1093));
  INV_X1    g0893(.A(G322), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n772), .A2(new_n778), .B1(new_n775), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1093), .B1(new_n603), .B2(new_n764), .C1(new_n1095), .C2(KEYINPUT115), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT115), .B2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n476), .B2(new_n768), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n767), .A2(new_n781), .B1(new_n761), .B2(new_n976), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1049), .A2(G303), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1086), .A2(new_n1092), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n751), .B1(new_n1083), .B2(new_n1084), .C1(new_n1103), .C2(new_n758), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n999), .B2(new_n807), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n745), .B1(new_n1077), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1075), .A2(KEYINPUT113), .A3(new_n1076), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1082), .A2(new_n1109), .ZN(G390));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n936), .B2(new_n911), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n930), .A2(new_n931), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n877), .B1(new_n721), .B2(new_n848), .ZN(new_n1114));
  OAI211_X1 g0914(.A(KEYINPUT117), .B(new_n912), .C1(new_n1114), .C2(new_n933), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n942), .A2(new_n737), .A3(G330), .A4(new_n738), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n678), .B1(new_n720), .B2(new_n710), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n877), .B1(new_n1120), .B2(new_n848), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n912), .B(new_n946), .C1(new_n1121), .C2(new_n933), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1116), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1119), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1113), .A2(new_n805), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n819), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n751), .B1(new_n1127), .B2(new_n256), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n776), .A2(G294), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n798), .A2(new_n830), .A3(new_n1129), .A4(new_n374), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n603), .A2(new_n781), .B1(new_n761), .B2(new_n778), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(G77), .C2(new_n765), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n220), .B2(new_n768), .C1(new_n426), .C2(new_n788), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT120), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n374), .B1(new_n776), .B2(G125), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1136), .B1(new_n228), .B2(new_n779), .C1(new_n761), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G132), .B2(new_n782), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1140));
  OR3_X1    g0940(.A1(new_n772), .A2(new_n1140), .A3(new_n835), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n772), .B2(new_n835), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n792), .C2(new_n764), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n796), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1139), .B(new_n1145), .C1(new_n960), .C2(new_n788), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1135), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1128), .B1(new_n1148), .B2(new_n757), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1125), .A2(new_n748), .B1(new_n1126), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n737), .A2(G330), .A3(new_n738), .A4(new_n848), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n933), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1152), .A2(new_n1117), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1114), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n868), .A3(new_n950), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1118), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1116), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n723), .A2(new_n449), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n669), .A3(new_n950), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1114), .B1(new_n1152), .B2(new_n1117), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1121), .B2(new_n1154), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1157), .A2(new_n1166), .A3(new_n702), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n1167), .ZN(G378));
  AND3_X1   g0968(.A1(new_n932), .A2(new_n938), .A3(KEYINPUT106), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT106), .B1(new_n932), .B2(new_n938), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT55), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n302), .B(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n270), .A2(new_n871), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT123), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1173), .B(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1169), .A2(new_n1170), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n925), .B2(new_n939), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n949), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n925), .A2(new_n939), .A3(new_n1176), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(G330), .A3(new_n1182), .A4(new_n948), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1183), .A3(new_n748), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n751), .B1(new_n1127), .B2(G50), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n533), .A2(G41), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G50), .B(new_n1186), .C1(new_n257), .C2(new_n452), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT121), .Z(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n761), .B2(new_n603), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G107), .B2(new_n782), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n799), .A2(G58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n776), .A2(G283), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1052), .A2(new_n1192), .A3(new_n1193), .A4(new_n965), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n431), .B2(new_n796), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1191), .B(new_n1195), .C1(new_n220), .C2(new_n788), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1188), .B1(new_n1189), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n773), .A2(new_n1144), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n835), .B2(new_n764), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n781), .A2(new_n1137), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G125), .C2(new_n762), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n960), .B2(new_n768), .C1(new_n831), .C2(new_n788), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n799), .A2(G159), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1197), .B1(new_n1189), .B2(new_n1196), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1208), .B2(new_n757), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1176), .B2(new_n806), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1184), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1162), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1166), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1180), .A4(new_n1183), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n702), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1212), .B1(new_n1216), .B2(new_n1218), .ZN(G375));
  AOI21_X1  g1019(.A(new_n1155), .B1(new_n868), .B2(new_n950), .ZN(new_n1220));
  OR3_X1    g1020(.A1(new_n1220), .A2(new_n1165), .A3(new_n1021), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n768), .A2(new_n835), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1192), .B1(new_n1137), .B2(new_n775), .C1(new_n792), .C2(new_n772), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n363), .B(new_n1223), .C1(G50), .C2(new_n765), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n831), .B2(new_n761), .C1(new_n960), .C2(new_n781), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1222), .B(new_n1225), .C1(new_n1049), .C2(new_n1144), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n788), .A2(new_n603), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n768), .A2(new_n426), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1054), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n773), .A2(G97), .B1(new_n776), .B2(G303), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n374), .A4(new_n959), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n778), .A2(new_n781), .B1(new_n761), .B2(new_n476), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1227), .A2(new_n1228), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n757), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n751), .B1(new_n1127), .B2(G68), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT124), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n933), .B2(new_n805), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1155), .B2(new_n748), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1221), .A2(new_n1239), .ZN(G381));
  OR3_X1    g1040(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G387), .A2(G381), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1109), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G375), .A2(G378), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .ZN(G407));
  AND2_X1   g1046(.A1(new_n1217), .A2(new_n702), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT57), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1162), .B1(new_n1125), .B2(new_n1165), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1211), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1254), .ZN(G409));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1251), .A2(new_n702), .A3(new_n1217), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1257), .B2(new_n1212), .ZN(new_n1258));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1184), .A2(new_n1167), .A3(new_n1150), .A4(new_n1210), .ZN(new_n1262));
  AND4_X1   g1062(.A1(new_n1020), .A2(new_n1215), .A3(new_n1183), .A4(new_n1180), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1256), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1211), .A2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1263), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1260), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1268), .B(KEYINPUT126), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1269));
  OAI211_X1 g1069(.A(KEYINPUT125), .B(new_n1156), .C1(new_n1220), .C2(KEYINPUT60), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1165), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n703), .B1(new_n1220), .B2(KEYINPUT60), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1239), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(G384), .A3(new_n1239), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(G2897), .A3(new_n1279), .A4(new_n1260), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(G2897), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1275), .A2(G384), .A3(new_n1239), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1275), .B2(new_n1239), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1265), .A2(new_n1269), .A3(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(G396), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G390), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1244), .A2(new_n1287), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1036), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1036), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1291), .A2(new_n1292), .A3(KEYINPUT61), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1294));
  NOR4_X1   g1094(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1264), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1264), .B1(G375), .B2(G378), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1286), .B(new_n1293), .C1(new_n1295), .C2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1285), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1305));
  NOR4_X1   g1105(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1264), .A4(new_n1294), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1303), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1300), .B1(new_n1307), .B2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1294), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1245), .B2(new_n1258), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G375), .A2(G378), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1254), .A2(new_n1315), .A3(new_n1312), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1308), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1317), .B(new_n1318), .ZN(G402));
endmodule


