//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n207), .B(new_n208), .C1(G1gat), .C2(new_n205), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT96), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n205), .A2(G1gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(KEYINPUT95), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n211), .B2(KEYINPUT95), .ZN(new_n213));
  OAI21_X1  g012(.A(G8gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT91), .B1(new_n217), .B2(new_n218), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT93), .ZN(new_n225));
  NOR3_X1   g024(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n229), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n231), .A2(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n221), .A2(new_n222), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G29gat), .A2(G36gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n227), .A2(KEYINPUT90), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n228), .B1(new_n226), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n223), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(KEYINPUT94), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT94), .B1(new_n233), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n216), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n240), .A3(new_n215), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n204), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n241), .A2(KEYINPUT17), .A3(new_n242), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT17), .A3(new_n239), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n216), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n202), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n240), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n216), .B(new_n250), .C1(new_n255), .C2(KEYINPUT17), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n247), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT89), .B(G197gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT11), .B(G169gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT12), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n254), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n254), .B2(new_n257), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT97), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n253), .ZN(new_n268));
  INV_X1    g067(.A(new_n248), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n257), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n263), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n257), .A3(new_n263), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT97), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n279), .A2(new_n280), .B1(G169gat), .B2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT66), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n291));
  INV_X1    g090(.A(new_n282), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n286), .A2(new_n287), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n280), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT67), .B1(new_n301), .B2(new_n302), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT28), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n300), .ZN(new_n325));
  AND2_X1   g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n278), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n324), .A2(KEYINPUT68), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT68), .B1(new_n324), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n314), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n277), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n312), .B1(new_n304), .B2(new_n305), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n330), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT68), .A3(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n338), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT75), .A3(new_n335), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n306), .A2(new_n313), .B1(new_n324), .B2(new_n330), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n335), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G197gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G197gat), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n354), .A2(new_n356), .A3(G204gat), .ZN(new_n357));
  AOI21_X1  g156(.A(G204gat), .B1(new_n354), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G211gat), .B(G218gat), .Z(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n360), .ZN(new_n362));
  INV_X1    g161(.A(G204gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n355), .A2(G197gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(new_n356), .A3(G204gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n368), .B2(new_n352), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n335), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n314), .A2(new_n333), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n372), .A2(KEYINPUT76), .B1(new_n336), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n370), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n335), .C1(new_n347), .C2(KEYINPUT29), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT77), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND4_X1  g181(.A1(new_n371), .A2(new_n378), .A3(KEYINPUT30), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n371), .B2(new_n378), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(new_n336), .ZN(new_n387));
  AND4_X1   g186(.A1(new_n375), .A2(new_n386), .A3(new_n377), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n345), .A2(new_n335), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n348), .B1(new_n389), .B2(new_n277), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n375), .B1(new_n390), .B2(new_n346), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT30), .A4(new_n382), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n276), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G134gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G127gat), .ZN(new_n403));
  INV_X1    g202(.A(G127gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G134gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT69), .ZN(new_n407));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(G113gat), .A2(G120gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(G113gat), .A2(G120gat), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT70), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT1), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n407), .A2(new_n410), .A3(new_n413), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n412), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n406), .B1(new_n420), .B2(KEYINPUT1), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G141gat), .B(G148gat), .Z(new_n423));
  INV_X1    g222(.A(G155gat), .ZN(new_n424));
  INV_X1    g223(.A(G162gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(KEYINPUT2), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G141gat), .B(G148gat), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n427), .B(new_n426), .C1(new_n431), .C2(KEYINPUT2), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n422), .B1(KEYINPUT3), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT80), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT80), .B1(new_n430), .B2(new_n432), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n419), .A2(new_n432), .A3(new_n430), .A4(new_n421), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n444), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n411), .A2(new_n415), .A3(new_n417), .A4(new_n412), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n409), .B2(new_n408), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n451), .B2(new_n407), .ZN(new_n452));
  INV_X1    g251(.A(new_n433), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(KEYINPUT83), .A3(new_n453), .A4(new_n446), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n448), .A2(new_n454), .A3(KEYINPUT84), .A4(new_n455), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n439), .B(new_n443), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n445), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n438), .B2(new_n422), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT5), .B1(new_n462), .B2(new_n440), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(KEYINPUT4), .A3(new_n453), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n446), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n440), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n439), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n433), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n435), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n422), .B(new_n470), .C1(new_n473), .C2(new_n469), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n441), .B1(new_n461), .B2(KEYINPUT4), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT82), .A4(new_n466), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n463), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n401), .B1(new_n460), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n468), .A2(new_n476), .ZN(new_n479));
  INV_X1    g278(.A(new_n463), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n459), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n474), .A3(new_n442), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n483), .A3(new_n400), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(KEYINPUT6), .B(new_n401), .C1(new_n460), .C2(new_n477), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n371), .A2(new_n378), .ZN(new_n490));
  INV_X1    g289(.A(new_n382), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n385), .A2(new_n394), .A3(new_n276), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n396), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n452), .B1(new_n339), .B2(new_n344), .ZN(new_n497));
  INV_X1    g296(.A(new_n303), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n293), .A2(new_n296), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(KEYINPUT66), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT25), .B1(new_n500), .B2(new_n298), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n333), .B(new_n422), .C1(new_n501), .C2(new_n312), .ZN(new_n502));
  INV_X1    g301(.A(G227gat), .ZN(new_n503));
  INV_X1    g302(.A(G233gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G15gat), .B(G43gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT71), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT33), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(KEYINPUT32), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n506), .A2(new_n514), .A3(KEYINPUT32), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g316(.A(new_n506), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n517), .B(new_n510), .C1(new_n518), .C2(KEYINPUT33), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT34), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n497), .A2(new_n502), .ZN(new_n522));
  INV_X1    g321(.A(new_n505), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT34), .B(new_n505), .C1(new_n497), .C2(new_n502), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(new_n526), .A3(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G78gat), .B(G106gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G228gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n338), .B1(new_n361), .B2(new_n369), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n473), .B1(new_n536), .B2(new_n469), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n338), .B1(new_n433), .B2(KEYINPUT3), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n370), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n370), .A2(new_n538), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT29), .B1(new_n369), .B2(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n359), .A2(new_n360), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n368), .A2(new_n362), .A3(new_n352), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT85), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT3), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n534), .B(new_n541), .C1(new_n547), .C2(new_n453), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n540), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n533), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n541), .A2(new_n534), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n542), .A2(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n469), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n433), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT29), .B1(new_n543), .B2(new_n544), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n438), .B1(new_n558), .B2(KEYINPUT3), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n534), .B1(new_n559), .B2(new_n541), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n549), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n532), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n530), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT35), .B1(new_n496), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n528), .B2(new_n529), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n529), .A2(new_n569), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT87), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n516), .A2(new_n526), .A3(new_n519), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n526), .B1(new_n516), .B2(new_n519), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT73), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n553), .A2(new_n563), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n486), .B2(new_n487), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n385), .A3(new_n394), .A4(new_n492), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n568), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  AOI211_X1 g384(.A(KEYINPUT88), .B(new_n583), .C1(new_n573), .C2(new_n578), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n567), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n576), .A2(new_n588), .A3(new_n571), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n488), .B1(new_n392), .B2(new_n382), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n375), .B1(new_n374), .B2(new_n377), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n593), .A2(KEYINPUT86), .B1(new_n370), .B2(new_n350), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n593), .A2(KEYINPUT86), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT37), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n382), .B1(new_n392), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT38), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n598), .A2(KEYINPUT38), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n592), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n462), .B2(new_n440), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n439), .B1(new_n458), .B2(new_n459), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n440), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n606), .A2(new_n400), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n605), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n607), .A2(KEYINPUT40), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT40), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  INV_X1    g409(.A(new_n478), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n385), .A2(new_n394), .A3(new_n492), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n564), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n591), .B1(new_n602), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n496), .A2(new_n564), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n275), .B1(new_n587), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G57gat), .B(G64gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT9), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G71gat), .ZN(new_n623));
  INV_X1    g422(.A(G78gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n621), .C1(KEYINPUT98), .C2(new_n620), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n622), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n622), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n622), .A2(new_n626), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n216), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n640), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G190gat), .B(G218gat), .Z(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(G85gat), .ZN(new_n654));
  INV_X1    g453(.A(G92gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n654), .A2(new_n655), .B1(KEYINPUT8), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  INV_X1    g457(.A(G85gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n655), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT7), .ZN(new_n661));
  NAND3_X1  g460(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(KEYINPUT7), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n657), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G99gat), .B(G106gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n657), .A2(new_n661), .A3(new_n665), .A4(new_n663), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n250), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n249), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n255), .B2(new_n669), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n653), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n241), .A2(new_n242), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n250), .B(new_n669), .C1(new_n255), .C2(KEYINPUT17), .ZN(new_n678));
  INV_X1    g477(.A(new_n653), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n652), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n674), .A2(new_n652), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(G230gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n504), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT104), .B(KEYINPUT10), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n629), .A2(new_n632), .A3(new_n669), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n676), .A2(new_n627), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n629), .A3(KEYINPUT10), .A4(new_n632), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n686), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(G120gat), .B(G148gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(G176gat), .B(G204gat), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n694), .A2(new_n696), .A3(new_n700), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n648), .A2(new_n684), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n707));
  INV_X1    g506(.A(new_n683), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n681), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n647), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n705), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n618), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n488), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT106), .B(G1gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1324gat));
  XOR2_X1   g516(.A(KEYINPUT16), .B(G8gat), .Z(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n618), .A2(new_n613), .A3(new_n713), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT108), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  INV_X1    g521(.A(new_n613), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n714), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n618), .A2(KEYINPUT107), .A3(new_n613), .A4(new_n713), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(G8gat), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n718), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n721), .B(new_n726), .C1(new_n728), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g528(.A(new_n591), .ZN(new_n730));
  OAI21_X1  g529(.A(G15gat), .B1(new_n714), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n579), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(G15gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n714), .B2(new_n733), .ZN(G1326gat));
  INV_X1    g533(.A(new_n564), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n714), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT43), .B(G22gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n684), .A2(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n385), .A2(new_n394), .A3(new_n276), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(new_n395), .A3(new_n493), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n580), .B1(new_n742), .B2(new_n565), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT87), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n577), .B1(new_n576), .B2(new_n571), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n584), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT88), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n579), .A2(new_n568), .A3(new_n584), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n615), .A2(new_n616), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n647), .A2(new_n705), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n264), .A2(new_n265), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT110), .B1(new_n742), .B2(new_n735), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n496), .A2(new_n756), .A3(new_n564), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n615), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n684), .B1(new_n587), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n751), .B(new_n754), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n488), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n752), .A2(new_n684), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n618), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n488), .A2(G29gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n618), .A2(new_n768), .A3(new_n762), .A4(new_n764), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(G1328gat));
  NOR3_X1   g571(.A1(new_n763), .A2(G36gat), .A3(new_n723), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g573(.A(G36gat), .B1(new_n760), .B2(new_n723), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1329gat));
  OAI21_X1  g575(.A(G43gat), .B1(new_n760), .B2(new_n730), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n763), .A2(G43gat), .A3(new_n732), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1330gat));
  NOR2_X1   g582(.A1(new_n763), .A2(new_n735), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n564), .A2(G50gat), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n784), .A2(G50gat), .B1(new_n760), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g586(.A1(new_n587), .A2(new_n758), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n710), .A2(new_n753), .A3(new_n704), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n488), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n789), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n723), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  AND2_X1   g595(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n795), .B2(new_n796), .ZN(G1333gat));
  NAND3_X1  g598(.A1(new_n790), .A2(new_n623), .A3(new_n579), .ZN(new_n800));
  OAI21_X1  g599(.A(G71gat), .B1(new_n794), .B2(new_n730), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g602(.A1(new_n794), .A2(new_n735), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(new_n624), .ZN(G1335gat));
  INV_X1    g604(.A(new_n753), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n648), .ZN(new_n807));
  AND4_X1   g606(.A1(KEYINPUT51), .A2(new_n788), .A3(new_n709), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n759), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT112), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n755), .A2(new_n615), .A3(new_n757), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n709), .B(new_n807), .C1(new_n811), .C2(new_n749), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n791), .A2(new_n654), .A3(new_n704), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n807), .A2(new_n704), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT111), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n751), .B(new_n820), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n488), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n817), .A2(new_n818), .B1(new_n654), .B2(new_n822), .ZN(G1336gat));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n788), .A2(new_n709), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n739), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n613), .A3(new_n751), .A4(new_n820), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n807), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n723), .A2(G92gat), .A3(new_n705), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n827), .A2(G92gat), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n830), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n810), .B2(new_n816), .ZN(new_n833));
  OAI21_X1  g632(.A(G92gat), .B1(new_n821), .B2(new_n723), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n824), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n824), .A2(new_n831), .B1(new_n833), .B2(new_n835), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n821), .B2(new_n730), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n732), .A2(G99gat), .A3(new_n705), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT113), .Z(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n817), .B2(new_n839), .ZN(G1338gat));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n564), .A3(new_n751), .A4(new_n820), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n705), .A2(new_n735), .A3(G106gat), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n842), .A2(G106gat), .B1(new_n829), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n843), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n810), .B2(new_n816), .ZN(new_n846));
  OAI21_X1  g645(.A(G106gat), .B1(new_n821), .B2(new_n735), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n841), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n841), .A2(new_n844), .B1(new_n846), .B2(new_n848), .ZN(G1339gat));
  OAI211_X1 g648(.A(new_n686), .B(new_n692), .C1(new_n695), .C2(new_n688), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n694), .A3(KEYINPUT54), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n852), .B(new_n687), .C1(new_n691), .C2(new_n693), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n701), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n703), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n701), .A3(new_n853), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n856), .B(new_n859), .C1(new_n264), .C2(new_n265), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n202), .B1(new_n256), .B2(new_n247), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n243), .A2(new_n247), .A3(new_n204), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n262), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n273), .A2(new_n704), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n709), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n855), .B1(new_n858), .B2(new_n857), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n273), .A2(new_n863), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n709), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n647), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n710), .A2(new_n753), .A3(new_n705), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n488), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n723), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n732), .A2(new_n564), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(G113gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n874), .A2(new_n875), .A3(new_n275), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n871), .A2(new_n723), .A3(new_n565), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n806), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n876), .A2(new_n879), .ZN(G1340gat));
  OR3_X1    g679(.A1(new_n877), .A2(G120gat), .A3(new_n705), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n871), .A2(new_n723), .A3(new_n704), .A4(new_n873), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n883), .A3(G120gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n882), .B2(G120gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT115), .Z(G1341gat));
  NOR3_X1   g686(.A1(new_n874), .A2(new_n404), .A3(new_n647), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n878), .A2(new_n648), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  AOI21_X1  g689(.A(G127gat), .B1(new_n889), .B2(KEYINPUT116), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1342gat));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n877), .A2(G134gat), .A3(new_n684), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n709), .A3(new_n873), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n893), .A2(new_n894), .B1(new_n895), .B2(G134gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n684), .A2(G134gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n872), .A2(new_n565), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT56), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n898), .B2(KEYINPUT56), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT118), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n896), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1343gat));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n871), .A2(new_n564), .A3(new_n730), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n723), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n275), .ZN(new_n914));
  INV_X1    g713(.A(G141gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n908), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n613), .A2(new_n488), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n730), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g718(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n869), .A2(new_n870), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n564), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n850), .A2(new_n694), .A3(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n853), .A2(new_n701), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n851), .A2(KEYINPUT120), .A3(new_n701), .A4(new_n853), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n858), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n856), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n266), .B1(new_n264), .B2(new_n265), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n272), .A2(KEYINPUT97), .A3(new_n273), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n864), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n684), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n868), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n648), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n870), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT57), .B(new_n564), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n919), .B1(new_n924), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n915), .B1(new_n941), .B2(new_n914), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n909), .A2(new_n613), .A3(new_n916), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n806), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(G141gat), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n917), .A2(new_n942), .B1(new_n945), .B2(new_n908), .ZN(G1344gat));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n735), .B(new_n920), .C1(new_n869), .C2(new_n870), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n707), .A2(new_n275), .A3(new_n712), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n564), .B1(new_n938), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT57), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n919), .A2(new_n705), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(G148gat), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n919), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n564), .A2(KEYINPUT57), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n930), .A2(new_n856), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n267), .B2(new_n274), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n709), .B1(new_n959), .B2(new_n864), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n647), .B1(new_n960), .B2(new_n868), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n870), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n704), .B(new_n956), .C1(new_n962), .C2(new_n923), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G148gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n955), .A2(KEYINPUT59), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n705), .A2(G148gat), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n911), .A2(new_n723), .A3(new_n912), .A4(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n947), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n948), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n707), .A2(new_n275), .A3(new_n712), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n735), .B1(new_n961), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n974), .B2(KEYINPUT57), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n953), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n964), .B1(new_n976), .B2(G148gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n965), .B1(new_n941), .B2(new_n704), .ZN(new_n978));
  OAI211_X1 g777(.A(KEYINPUT122), .B(new_n969), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n971), .A2(new_n979), .ZN(G1345gat));
  NAND4_X1  g779(.A1(new_n911), .A2(new_n723), .A3(new_n648), .A4(new_n912), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(G155gat), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n647), .A2(new_n424), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n941), .B2(new_n985), .ZN(G1346gat));
  INV_X1    g785(.A(new_n913), .ZN(new_n987));
  AOI21_X1  g786(.A(G162gat), .B1(new_n987), .B2(new_n709), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n684), .A2(new_n425), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n941), .B2(new_n989), .ZN(G1347gat));
  NOR2_X1   g789(.A1(new_n723), .A2(new_n791), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n922), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n992), .A2(new_n565), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(new_n294), .A3(new_n806), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n873), .ZN(new_n995));
  OAI21_X1  g794(.A(G169gat), .B1(new_n995), .B2(new_n275), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1348gat));
  NAND3_X1  g796(.A1(new_n993), .A2(new_n284), .A3(new_n704), .ZN(new_n998));
  OAI21_X1  g797(.A(G176gat), .B1(new_n995), .B2(new_n705), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1349gat));
  NAND4_X1  g799(.A1(new_n993), .A2(new_n316), .A3(new_n318), .A4(new_n648), .ZN(new_n1001));
  OAI21_X1  g800(.A(G183gat), .B1(new_n995), .B2(new_n647), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT124), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g803(.A1(new_n993), .A2(new_n319), .A3(new_n709), .ZN(new_n1005));
  OAI21_X1  g804(.A(G190gat), .B1(new_n995), .B2(new_n684), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1351gat));
  NAND2_X1  g808(.A1(new_n730), .A2(new_n991), .ZN(new_n1010));
  INV_X1    g809(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n922), .A2(new_n564), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g811(.A(G197gat), .B1(new_n1012), .B2(new_n806), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n952), .A2(new_n1010), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n275), .A2(new_n353), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(G1352gat));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n704), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1014), .A2(KEYINPUT126), .A3(new_n704), .ZN(new_n1020));
  XOR2_X1   g819(.A(KEYINPUT125), .B(G204gat), .Z(new_n1021));
  NAND3_X1  g820(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n705), .A2(new_n1021), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1012), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g823(.A(new_n1024), .B(KEYINPUT62), .Z(new_n1025));
  NAND2_X1  g824(.A1(new_n1022), .A2(new_n1025), .ZN(G1353gat));
  INV_X1    g825(.A(G211gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n1027), .A3(new_n648), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1014), .A2(new_n648), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  AND2_X1   g831(.A1(new_n1014), .A2(KEYINPUT127), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n709), .B1(new_n1014), .B2(KEYINPUT127), .ZN(new_n1034));
  OAI21_X1  g833(.A(G218gat), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g834(.A(G218gat), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n1012), .A2(new_n1036), .A3(new_n709), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1035), .A2(new_n1037), .ZN(G1355gat));
endmodule


