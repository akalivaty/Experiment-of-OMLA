

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752;

  XOR2_X1 U365 ( .A(KEYINPUT124), .B(n715), .Z(n716) );
  NOR2_X1 U366 ( .A1(n374), .A2(n542), .ZN(n346) );
  NAND2_X2 U367 ( .A1(n405), .A2(n547), .ZN(n548) );
  NOR2_X2 U368 ( .A1(n750), .A2(n345), .ZN(n582) );
  INV_X1 U369 ( .A(n580), .ZN(n345) );
  XNOR2_X2 U370 ( .A(n539), .B(n538), .ZN(n580) );
  XNOR2_X2 U371 ( .A(n579), .B(n578), .ZN(n750) );
  NAND2_X1 U372 ( .A1(n346), .A2(n485), .ZN(n486) );
  XNOR2_X1 U373 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n376) );
  INV_X1 U374 ( .A(n641), .ZN(n638) );
  AND2_X2 U375 ( .A1(n384), .A2(n382), .ZN(n381) );
  XNOR2_X2 U376 ( .A(n548), .B(KEYINPUT108), .ZN(n563) );
  XNOR2_X2 U377 ( .A(n434), .B(n370), .ZN(n674) );
  NOR2_X1 U378 ( .A1(n639), .A2(n678), .ZN(n390) );
  AND2_X1 U379 ( .A1(n392), .A2(n649), .ZN(n391) );
  XNOR2_X1 U380 ( .A(n413), .B(n574), .ZN(n749) );
  XNOR2_X1 U381 ( .A(n554), .B(n553), .ZN(n645) );
  AND2_X1 U382 ( .A1(n551), .A2(n398), .ZN(n670) );
  NOR2_X1 U383 ( .A1(n677), .A2(n676), .ZN(n367) );
  XNOR2_X1 U384 ( .A(n393), .B(n737), .ZN(n719) );
  XNOR2_X1 U385 ( .A(n594), .B(KEYINPUT86), .ZN(n595) );
  INV_X1 U386 ( .A(KEYINPUT41), .ZN(n366) );
  OR2_X1 U387 ( .A1(n558), .A2(n529), .ZN(n676) );
  BUF_X1 U388 ( .A(n704), .Z(n347) );
  NOR2_X2 U389 ( .A1(n549), .A2(n532), .ZN(n417) );
  NOR2_X2 U390 ( .A1(n549), .A2(n532), .ZN(n356) );
  XNOR2_X2 U391 ( .A(n528), .B(KEYINPUT0), .ZN(n549) );
  XNOR2_X1 U392 ( .A(n455), .B(n454), .ZN(n478) );
  XNOR2_X1 U393 ( .A(G128), .B(G119), .ZN(n440) );
  XOR2_X1 U394 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n444) );
  XNOR2_X1 U395 ( .A(n414), .B(G110), .ZN(n457) );
  INV_X1 U396 ( .A(G107), .ZN(n414) );
  INV_X1 U397 ( .A(n673), .ZN(n402) );
  NOR2_X1 U398 ( .A1(n575), .A2(n542), .ZN(n587) );
  XNOR2_X1 U399 ( .A(n481), .B(n480), .ZN(n588) );
  NOR2_X2 U400 ( .A1(n719), .A2(G902), .ZN(n451) );
  INV_X1 U401 ( .A(n659), .ZN(n404) );
  INV_X1 U402 ( .A(n541), .ZN(n575) );
  AND2_X1 U403 ( .A1(n359), .A2(n659), .ZN(n577) );
  BUF_X2 U404 ( .A(n588), .Z(n398) );
  XNOR2_X1 U405 ( .A(G140), .B(G104), .ZN(n462) );
  XNOR2_X1 U406 ( .A(n390), .B(KEYINPUT47), .ZN(n389) );
  INV_X1 U407 ( .A(KEYINPUT44), .ZN(n364) );
  XNOR2_X1 U408 ( .A(G137), .B(KEYINPUT76), .ZN(n471) );
  XOR2_X1 U409 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n472) );
  XNOR2_X1 U410 ( .A(G119), .B(KEYINPUT3), .ZN(n426) );
  INV_X1 U411 ( .A(KEYINPUT77), .ZN(n373) );
  NAND2_X1 U412 ( .A1(n432), .A2(KEYINPUT2), .ZN(n386) );
  XOR2_X1 U413 ( .A(G131), .B(G134), .Z(n738) );
  XOR2_X1 U414 ( .A(G137), .B(KEYINPUT70), .Z(n456) );
  XNOR2_X1 U415 ( .A(n453), .B(G125), .ZN(n438) );
  XOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n422) );
  NOR2_X1 U417 ( .A1(n667), .A2(n398), .ZN(n668) );
  INV_X1 U418 ( .A(KEYINPUT38), .ZN(n370) );
  XNOR2_X1 U419 ( .A(n483), .B(KEYINPUT30), .ZN(n374) );
  INV_X1 U420 ( .A(G902), .ZN(n499) );
  XNOR2_X1 U421 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U422 ( .A(n442), .B(n445), .ZN(n394) );
  INV_X1 U423 ( .A(G128), .ZN(n418) );
  XNOR2_X1 U424 ( .A(G134), .B(G116), .ZN(n487) );
  XOR2_X1 U425 ( .A(G107), .B(G122), .Z(n488) );
  XNOR2_X1 U426 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n489) );
  XOR2_X1 U427 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n490) );
  XOR2_X1 U428 ( .A(G104), .B(G122), .Z(n507) );
  XNOR2_X1 U429 ( .A(n416), .B(n438), .ZN(n506) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n416) );
  INV_X1 U431 ( .A(G140), .ZN(n375) );
  XNOR2_X1 U432 ( .A(G143), .B(G131), .ZN(n503) );
  XOR2_X1 U433 ( .A(KEYINPUT100), .B(G113), .Z(n504) );
  XNOR2_X1 U434 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U435 ( .A(n457), .ZN(n458) );
  NOR2_X1 U436 ( .A1(n565), .A2(n566), .ZN(n570) );
  NAND2_X1 U437 ( .A1(n380), .A2(n379), .ZN(n378) );
  NOR2_X1 U438 ( .A1(n663), .A2(n402), .ZN(n401) );
  INV_X1 U439 ( .A(KEYINPUT36), .ZN(n594) );
  NAND2_X1 U440 ( .A1(n412), .A2(n409), .ZN(n411) );
  XNOR2_X1 U441 ( .A(n396), .B(KEYINPUT28), .ZN(n590) );
  NAND2_X1 U442 ( .A1(n587), .A2(n397), .ZN(n396) );
  AND2_X1 U443 ( .A1(n398), .A2(n530), .ZN(n397) );
  NOR2_X1 U444 ( .A1(n404), .A2(n543), .ZN(n403) );
  NOR2_X1 U445 ( .A1(n575), .A2(n398), .ZN(n576) );
  INV_X1 U446 ( .A(n398), .ZN(n556) );
  XNOR2_X1 U447 ( .A(n347), .B(n703), .ZN(n705) );
  AND2_X1 U448 ( .A1(n613), .A2(n615), .ZN(n348) );
  NOR2_X1 U449 ( .A1(n412), .A2(n557), .ZN(n349) );
  XNOR2_X1 U450 ( .A(n398), .B(KEYINPUT6), .ZN(n566) );
  AND2_X1 U451 ( .A1(n411), .A2(n573), .ZN(n350) );
  NAND2_X1 U452 ( .A1(n571), .A2(n572), .ZN(n351) );
  INV_X1 U453 ( .A(G146), .ZN(n453) );
  INV_X1 U454 ( .A(n572), .ZN(n409) );
  XNOR2_X1 U455 ( .A(n506), .B(n439), .ZN(n737) );
  XOR2_X1 U456 ( .A(n699), .B(n698), .Z(n352) );
  INV_X1 U457 ( .A(KEYINPUT78), .ZN(n615) );
  XNOR2_X1 U458 ( .A(G902), .B(KEYINPUT15), .ZN(n620) );
  XOR2_X1 U459 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n353) );
  OR2_X1 U460 ( .A1(n742), .A2(G952), .ZN(n700) );
  XNOR2_X1 U461 ( .A(n354), .B(n355), .ZN(n600) );
  NOR2_X1 U462 ( .A1(n699), .A2(n432), .ZN(n354) );
  NAND2_X1 U463 ( .A1(n482), .A2(G210), .ZN(n355) );
  BUF_X1 U464 ( .A(n701), .Z(n702) );
  XNOR2_X1 U465 ( .A(n367), .B(n366), .ZN(n689) );
  XOR2_X1 U466 ( .A(n709), .B(KEYINPUT59), .Z(n710) );
  XNOR2_X1 U467 ( .A(n603), .B(KEYINPUT40), .ZN(n415) );
  NAND2_X1 U468 ( .A1(n600), .A2(n673), .ZN(n521) );
  XNOR2_X1 U469 ( .A(n365), .B(n364), .ZN(n583) );
  NOR2_X1 U470 ( .A1(n619), .A2(n617), .ZN(n357) );
  BUF_X1 U471 ( .A(n415), .Z(n358) );
  XNOR2_X1 U472 ( .A(n356), .B(KEYINPUT22), .ZN(n359) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT22), .ZN(n546) );
  XNOR2_X1 U474 ( .A(n589), .B(n534), .ZN(n597) );
  NAND2_X1 U475 ( .A1(n597), .A2(n550), .ZN(n565) );
  NAND2_X1 U476 ( .A1(n381), .A2(n378), .ZN(n360) );
  NAND2_X1 U477 ( .A1(n381), .A2(n378), .ZN(n657) );
  BUF_X2 U478 ( .A(n600), .Z(n434) );
  NAND2_X1 U479 ( .A1(n701), .A2(G210), .ZN(n363) );
  XNOR2_X1 U480 ( .A(n361), .B(n353), .ZN(G51) );
  NAND2_X1 U481 ( .A1(n362), .A2(n700), .ZN(n361) );
  XNOR2_X1 U482 ( .A(n363), .B(n352), .ZN(n362) );
  XNOR2_X1 U483 ( .A(n406), .B(KEYINPUT85), .ZN(n405) );
  NAND2_X1 U484 ( .A1(n657), .A2(n387), .ZN(n621) );
  NAND2_X1 U485 ( .A1(n563), .A2(n368), .ZN(n564) );
  NAND2_X1 U486 ( .A1(n407), .A2(n350), .ZN(n413) );
  NAND2_X1 U487 ( .A1(n582), .A2(n749), .ZN(n365) );
  NAND2_X1 U488 ( .A1(n562), .A2(n561), .ZN(n368) );
  OR2_X2 U489 ( .A1(n412), .A2(n552), .ZN(n554) );
  NAND2_X1 U490 ( .A1(n415), .A2(n752), .ZN(n369) );
  XNOR2_X1 U491 ( .A(n369), .B(n607), .ZN(n371) );
  NOR2_X2 U492 ( .A1(n619), .A2(n617), .ZN(n614) );
  INV_X1 U493 ( .A(n571), .ZN(n412) );
  NAND2_X1 U494 ( .A1(n371), .A2(n608), .ZN(n609) );
  NAND2_X1 U495 ( .A1(n377), .A2(n372), .ZN(n385) );
  XNOR2_X1 U496 ( .A(n653), .B(n373), .ZN(n372) );
  NOR2_X1 U497 ( .A1(n651), .A2(n620), .ZN(n377) );
  AND2_X1 U498 ( .A1(n357), .A2(n348), .ZN(n379) );
  INV_X1 U499 ( .A(n651), .ZN(n380) );
  NAND2_X1 U500 ( .A1(n383), .A2(KEYINPUT78), .ZN(n382) );
  NAND2_X1 U501 ( .A1(n614), .A2(n613), .ZN(n383) );
  NAND2_X1 U502 ( .A1(n651), .A2(KEYINPUT78), .ZN(n384) );
  NAND2_X1 U503 ( .A1(n385), .A2(n386), .ZN(n387) );
  INV_X1 U504 ( .A(KEYINPUT2), .ZN(n388) );
  NAND2_X1 U505 ( .A1(n391), .A2(n389), .ZN(n599) );
  INV_X1 U506 ( .A(n592), .ZN(n392) );
  NAND2_X1 U507 ( .A1(n493), .A2(G221), .ZN(n395) );
  NOR2_X2 U508 ( .A1(n619), .A2(n618), .ZN(n653) );
  AND2_X1 U509 ( .A1(n543), .A2(n399), .ZN(n593) );
  NOR2_X1 U510 ( .A1(n638), .A2(n400), .ZN(n399) );
  NAND2_X1 U511 ( .A1(n587), .A2(n401), .ZN(n400) );
  NAND2_X1 U512 ( .A1(n546), .A2(n403), .ZN(n406) );
  OR2_X1 U513 ( .A1(n688), .A2(n409), .ZN(n408) );
  NAND2_X1 U514 ( .A1(n410), .A2(n408), .ZN(n407) );
  NAND2_X1 U515 ( .A1(n688), .A2(n351), .ZN(n410) );
  XNOR2_X2 U516 ( .A(n466), .B(n465), .ZN(n589) );
  XNOR2_X1 U517 ( .A(n358), .B(G131), .ZN(G33) );
  XNOR2_X2 U518 ( .A(n609), .B(KEYINPUT48), .ZN(n619) );
  NOR2_X2 U519 ( .A1(n712), .A2(n723), .ZN(n713) );
  INV_X1 U520 ( .A(n541), .ZN(n452) );
  XNOR2_X1 U521 ( .A(n431), .B(n731), .ZN(n699) );
  XNOR2_X1 U522 ( .A(n455), .B(n425), .ZN(n431) );
  INV_X1 U523 ( .A(KEYINPUT46), .ZN(n607) );
  INV_X1 U524 ( .A(n456), .ZN(n439) );
  XNOR2_X1 U525 ( .A(n479), .B(n622), .ZN(n480) );
  XNOR2_X1 U526 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n570), .B(n569), .ZN(n688) );
  BUF_X1 U528 ( .A(n651), .Z(n727) );
  BUF_X1 U529 ( .A(n653), .Z(n741) );
  INV_X1 U530 ( .A(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U531 ( .A(n596), .B(n595), .ZN(n598) );
  XNOR2_X1 U532 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X2 U533 ( .A(G143), .B(KEYINPUT65), .ZN(n419) );
  XNOR2_X2 U534 ( .A(n419), .B(n418), .ZN(n496) );
  XNOR2_X2 U535 ( .A(n496), .B(KEYINPUT4), .ZN(n739) );
  XNOR2_X2 U536 ( .A(n739), .B(G101), .ZN(n455) );
  INV_X1 U537 ( .A(KEYINPUT64), .ZN(n420) );
  XNOR2_X2 U538 ( .A(n420), .B(G953), .ZN(n742) );
  NAND2_X1 U539 ( .A1(n742), .A2(G224), .ZN(n421) );
  XNOR2_X1 U540 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U541 ( .A(n438), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U542 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U543 ( .A(G113), .B(G116), .Z(n427) );
  XNOR2_X1 U544 ( .A(n427), .B(n426), .ZN(n474) );
  INV_X1 U545 ( .A(n507), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n474), .B(n428), .ZN(n430) );
  XNOR2_X1 U547 ( .A(n457), .B(KEYINPUT16), .ZN(n429) );
  XNOR2_X1 U548 ( .A(n430), .B(n429), .ZN(n731) );
  INV_X1 U549 ( .A(n620), .ZN(n432) );
  INV_X1 U550 ( .A(G237), .ZN(n433) );
  NAND2_X1 U551 ( .A1(n499), .A2(n433), .ZN(n482) );
  INV_X1 U552 ( .A(n434), .ZN(n520) );
  NAND2_X1 U553 ( .A1(G234), .A2(n620), .ZN(n435) );
  XNOR2_X1 U554 ( .A(KEYINPUT20), .B(n435), .ZN(n446) );
  AND2_X1 U555 ( .A1(n446), .A2(G221), .ZN(n437) );
  XNOR2_X1 U556 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n436) );
  XNOR2_X1 U557 ( .A(n437), .B(n436), .ZN(n663) );
  INV_X1 U558 ( .A(n663), .ZN(n530) );
  XOR2_X1 U559 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n441) );
  XNOR2_X1 U560 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U561 ( .A(G110), .B(KEYINPUT23), .Z(n445) );
  NAND2_X1 U562 ( .A1(G234), .A2(n742), .ZN(n443) );
  XNOR2_X1 U563 ( .A(n444), .B(n443), .ZN(n493) );
  XOR2_X1 U564 ( .A(KEYINPUT94), .B(KEYINPUT80), .Z(n448) );
  NAND2_X1 U565 ( .A1(n446), .A2(G217), .ZN(n447) );
  XNOR2_X1 U566 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U567 ( .A(KEYINPUT25), .B(n449), .ZN(n450) );
  XNOR2_X2 U568 ( .A(n451), .B(n450), .ZN(n541) );
  NAND2_X1 U569 ( .A1(n530), .A2(n452), .ZN(n658) );
  XOR2_X1 U570 ( .A(G146), .B(n738), .Z(n454) );
  XOR2_X1 U571 ( .A(n456), .B(KEYINPUT81), .Z(n461) );
  NAND2_X1 U572 ( .A1(G227), .A2(n742), .ZN(n459) );
  XNOR2_X1 U573 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U574 ( .A(n478), .B(n464), .ZN(n704) );
  OR2_X2 U575 ( .A1(n704), .A2(G902), .ZN(n466) );
  XOR2_X1 U576 ( .A(KEYINPUT72), .B(G469), .Z(n465) );
  NOR2_X2 U577 ( .A1(n658), .A2(n589), .ZN(n555) );
  XNOR2_X1 U578 ( .A(n555), .B(KEYINPUT112), .ZN(n485) );
  NAND2_X1 U579 ( .A1(G234), .A2(G237), .ZN(n467) );
  XNOR2_X1 U580 ( .A(n467), .B(KEYINPUT14), .ZN(n468) );
  NAND2_X1 U581 ( .A1(G952), .A2(n468), .ZN(n687) );
  NOR2_X1 U582 ( .A1(G953), .A2(n687), .ZN(n525) );
  NAND2_X1 U583 ( .A1(G902), .A2(n468), .ZN(n523) );
  OR2_X1 U584 ( .A1(n742), .A2(n523), .ZN(n469) );
  NOR2_X1 U585 ( .A1(G900), .A2(n469), .ZN(n470) );
  NOR2_X1 U586 ( .A1(n525), .A2(n470), .ZN(n542) );
  XNOR2_X1 U587 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U588 ( .A(n474), .B(n473), .Z(n476) );
  NOR2_X1 U589 ( .A1(G953), .A2(G237), .ZN(n508) );
  NAND2_X1 U590 ( .A1(n508), .A2(G210), .ZN(n475) );
  XOR2_X1 U591 ( .A(n476), .B(n475), .Z(n477) );
  XNOR2_X1 U592 ( .A(n478), .B(n477), .ZN(n623) );
  NOR2_X1 U593 ( .A1(n623), .A2(G902), .ZN(n481) );
  XNOR2_X1 U594 ( .A(KEYINPUT75), .B(KEYINPUT97), .ZN(n479) );
  INV_X1 U595 ( .A(G472), .ZN(n622) );
  NAND2_X1 U596 ( .A1(n482), .A2(G214), .ZN(n673) );
  NAND2_X1 U597 ( .A1(n588), .A2(n673), .ZN(n483) );
  XNOR2_X2 U598 ( .A(n486), .B(KEYINPUT79), .ZN(n601) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U600 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U601 ( .A(n492), .B(n491), .Z(n495) );
  NAND2_X1 U602 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n498) );
  INV_X1 U604 ( .A(n496), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n498), .B(n497), .ZN(n715) );
  NAND2_X1 U606 ( .A1(n715), .A2(n499), .ZN(n502) );
  INV_X1 U607 ( .A(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U608 ( .A(n500), .B(G478), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n502), .B(n501), .ZN(n559) );
  INV_X1 U610 ( .A(n559), .ZN(n529) );
  XNOR2_X1 U611 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n516) );
  XNOR2_X1 U612 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U613 ( .A(n506), .B(n505), .ZN(n514) );
  XNOR2_X1 U614 ( .A(n507), .B(KEYINPUT99), .ZN(n512) );
  XOR2_X1 U615 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n510) );
  NAND2_X1 U616 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U617 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U618 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U619 ( .A(n514), .B(n513), .ZN(n709) );
  NOR2_X1 U620 ( .A1(G902), .A2(n709), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n518) );
  INV_X1 U622 ( .A(G475), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n558) );
  AND2_X1 U624 ( .A1(n529), .A2(n558), .ZN(n573) );
  NAND2_X1 U625 ( .A1(n601), .A2(n573), .ZN(n519) );
  NOR2_X1 U626 ( .A1(n520), .A2(n519), .ZN(n592) );
  XOR2_X1 U627 ( .A(G143), .B(n592), .Z(G45) );
  XNOR2_X2 U628 ( .A(n521), .B(KEYINPUT19), .ZN(n591) );
  XOR2_X1 U629 ( .A(G898), .B(KEYINPUT90), .Z(n726) );
  NAND2_X1 U630 ( .A1(n726), .A2(G953), .ZN(n522) );
  XOR2_X1 U631 ( .A(KEYINPUT91), .B(n522), .Z(n733) );
  NOR2_X1 U632 ( .A1(n523), .A2(n733), .ZN(n524) );
  OR2_X1 U633 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U634 ( .A(n526), .B(KEYINPUT92), .ZN(n527) );
  NAND2_X1 U635 ( .A1(n591), .A2(n527), .ZN(n528) );
  INV_X1 U636 ( .A(n676), .ZN(n531) );
  NAND2_X1 U637 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U638 ( .A(KEYINPUT107), .ZN(n533) );
  XNOR2_X1 U639 ( .A(n541), .B(n533), .ZN(n662) );
  NAND2_X1 U640 ( .A1(n566), .A2(n662), .ZN(n535) );
  INV_X1 U641 ( .A(n597), .ZN(n659) );
  NOR2_X1 U642 ( .A1(n535), .A2(n659), .ZN(n536) );
  NAND2_X1 U643 ( .A1(n359), .A2(n536), .ZN(n539) );
  INV_X1 U644 ( .A(KEYINPUT67), .ZN(n537) );
  XNOR2_X1 U645 ( .A(n537), .B(KEYINPUT32), .ZN(n538) );
  XNOR2_X1 U646 ( .A(n580), .B(G119), .ZN(G21) );
  NAND2_X1 U647 ( .A1(n559), .A2(n558), .ZN(n540) );
  XNOR2_X2 U648 ( .A(n540), .B(KEYINPUT105), .ZN(n641) );
  INV_X1 U649 ( .A(n566), .ZN(n543) );
  NAND2_X1 U650 ( .A1(n593), .A2(n659), .ZN(n544) );
  XOR2_X1 U651 ( .A(KEYINPUT43), .B(n544), .Z(n545) );
  NOR2_X1 U652 ( .A1(n545), .A2(n434), .ZN(n617) );
  XOR2_X1 U653 ( .A(n617), .B(G140), .Z(G42) );
  INV_X1 U654 ( .A(n662), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n563), .B(G101), .ZN(G3) );
  INV_X1 U656 ( .A(n658), .ZN(n550) );
  INV_X1 U657 ( .A(n565), .ZN(n551) );
  INV_X1 U658 ( .A(n670), .ZN(n552) );
  XNOR2_X1 U659 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n553) );
  NAND2_X1 U660 ( .A1(n556), .A2(n555), .ZN(n557) );
  OR2_X1 U661 ( .A1(n645), .A2(n349), .ZN(n562) );
  NOR2_X1 U662 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U663 ( .A(n560), .B(KEYINPUT106), .ZN(n644) );
  NOR2_X1 U664 ( .A1(n644), .A2(n641), .ZN(n678) );
  INV_X1 U665 ( .A(n678), .ZN(n561) );
  XNOR2_X1 U666 ( .A(n564), .B(KEYINPUT109), .ZN(n584) );
  XNOR2_X1 U667 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n567) );
  XNOR2_X1 U668 ( .A(n567), .B(KEYINPUT87), .ZN(n568) );
  XNOR2_X1 U669 ( .A(KEYINPUT111), .B(n568), .ZN(n569) );
  INV_X1 U670 ( .A(n549), .ZN(n571) );
  XOR2_X1 U671 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n572) );
  INV_X1 U672 ( .A(KEYINPUT35), .ZN(n574) );
  NAND2_X1 U673 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U674 ( .A(KEYINPUT110), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U676 ( .A(KEYINPUT45), .ZN(n585) );
  XNOR2_X2 U677 ( .A(n586), .B(n585), .ZN(n651) );
  NOR2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n604), .A2(n591), .ZN(n639) );
  NAND2_X1 U680 ( .A1(n593), .A2(n434), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n598), .A2(n404), .ZN(n649) );
  XNOR2_X1 U682 ( .A(n599), .B(KEYINPUT71), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n601), .A2(n674), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n602), .B(KEYINPUT39), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n610), .A2(n641), .ZN(n603) );
  XOR2_X1 U686 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n606) );
  NAND2_X1 U687 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U688 ( .A1(n604), .A2(n689), .ZN(n605) );
  XNOR2_X1 U689 ( .A(n606), .B(n605), .ZN(n752) );
  BUF_X1 U690 ( .A(n610), .Z(n611) );
  NAND2_X1 U691 ( .A1(n611), .A2(n644), .ZN(n650) );
  NAND2_X1 U692 ( .A1(n650), .A2(KEYINPUT2), .ZN(n612) );
  XOR2_X1 U693 ( .A(KEYINPUT82), .B(n612), .Z(n613) );
  INV_X1 U694 ( .A(n650), .ZN(n616) );
  OR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X2 U696 ( .A(n621), .B(KEYINPUT66), .ZN(n708) );
  NOR2_X1 U697 ( .A1(n708), .A2(n622), .ZN(n626) );
  XOR2_X1 U698 ( .A(KEYINPUT89), .B(KEYINPUT62), .Z(n624) );
  XNOR2_X1 U699 ( .A(n623), .B(n624), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n627), .A2(n700), .ZN(n629) );
  XNOR2_X1 U702 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(G57) );
  NAND2_X1 U704 ( .A1(n349), .A2(n641), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U707 ( .A1(n349), .A2(n644), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(G107), .B(n633), .ZN(G9) );
  INV_X1 U710 ( .A(n644), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n639), .A2(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT116), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(G128), .B(n637), .ZN(G30) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U716 ( .A(G146), .B(n640), .Z(G48) );
  XOR2_X1 U717 ( .A(G113), .B(KEYINPUT117), .Z(n643) );
  NAND2_X1 U718 ( .A1(n641), .A2(n645), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n646), .B(KEYINPUT118), .ZN(n647) );
  XNOR2_X1 U722 ( .A(G116), .B(n647), .ZN(G18) );
  XOR2_X1 U723 ( .A(G125), .B(KEYINPUT37), .Z(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(G27) );
  XNOR2_X1 U725 ( .A(G134), .B(n650), .ZN(G36) );
  XNOR2_X1 U726 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n697) );
  NAND2_X1 U727 ( .A1(n727), .A2(n388), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(KEYINPUT83), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n741), .A2(KEYINPUT2), .ZN(n654) );
  NOR2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n360), .A2(n656), .ZN(n695) );
  XOR2_X1 U732 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n661) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(n664), .Z(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(KEYINPUT120), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT51), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n672), .A2(n689), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT121), .B(n681), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n682), .A2(n688), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U749 ( .A(KEYINPUT52), .B(n685), .Z(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n691) );
  AND2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U753 ( .A(KEYINPUT122), .B(n692), .Z(n693) );
  NOR2_X1 U754 ( .A1(G953), .A2(n693), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(G75) );
  INV_X1 U757 ( .A(n708), .ZN(n701) );
  XOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n698) );
  INV_X1 U759 ( .A(n700), .ZN(n723) );
  NAND2_X1 U760 ( .A1(n702), .A2(G469), .ZN(n706) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  NOR2_X1 U762 ( .A1(n707), .A2(n723), .ZN(G54) );
  INV_X1 U763 ( .A(n708), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n714), .A2(G475), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n713), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U767 ( .A1(n702), .A2(G478), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n723), .A2(n718), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n702), .A2(G217), .ZN(n721) );
  XOR2_X1 U771 ( .A(n719), .B(KEYINPUT125), .Z(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(G66) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n724) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n724), .Z(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U777 ( .A1(n727), .A2(G953), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  NOR2_X1 U779 ( .A1(n730), .A2(n729), .ZN(n736) );
  XNOR2_X1 U780 ( .A(G101), .B(n731), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n732), .B(KEYINPUT127), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n736), .B(n735), .ZN(G69) );
  XOR2_X1 U784 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U785 ( .A(n737), .B(n740), .ZN(n744) );
  XOR2_X1 U786 ( .A(n744), .B(n741), .Z(n743) );
  NAND2_X1 U787 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U788 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U789 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U790 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U791 ( .A1(n748), .A2(n747), .ZN(G72) );
  XNOR2_X1 U792 ( .A(G122), .B(n749), .ZN(G24) );
  XNOR2_X1 U793 ( .A(G110), .B(KEYINPUT115), .ZN(n751) );
  XNOR2_X1 U794 ( .A(n751), .B(n750), .ZN(G12) );
  XNOR2_X1 U795 ( .A(G137), .B(n752), .ZN(G39) );
endmodule

