//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n472), .A2(KEYINPUT70), .A3(G137), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n469), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(G2105), .B2(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(new_n472), .B(KEYINPUT71), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT72), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n482), .A2(new_n469), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n466), .B2(new_n467), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(new_n504), .C1(new_n467), .C2(new_n466), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT73), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G543), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT74), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n513), .A2(new_n519), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n518), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n512), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n507), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n536), .B1(new_n511), .B2(new_n537), .C1(new_n538), .C2(new_n517), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(G43), .A2(new_n512), .B1(new_n518), .B2(G81), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n516), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n507), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(new_n546), .B2(new_n545), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n507), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n517), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n512), .A2(new_n561), .A3(G53), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n511), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  XNOR2_X1  g141(.A(new_n539), .B(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G301));
  NAND2_X1  g143(.A1(new_n512), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n518), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n512), .A2(G48), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G86), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n507), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n518), .A2(G85), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n512), .A2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n507), .C2(new_n580), .ZN(G290));
  NAND3_X1  g156(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n517), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n516), .A2(G66), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n512), .A2(G54), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT78), .B1(new_n592), .B2(G868), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n567), .A2(new_n594), .ZN(new_n595));
  MUX2_X1   g170(.A(new_n593), .B(KEYINPUT78), .S(new_n595), .Z(G284));
  MUX2_X1   g171(.A(new_n593), .B(KEYINPUT78), .S(new_n595), .Z(G321));
  NOR2_X1   g172(.A1(G286), .A2(new_n594), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n565), .B(KEYINPUT80), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n594), .ZN(G297));
  AOI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n594), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G860), .ZN(G148));
  OAI21_X1  g178(.A(KEYINPUT81), .B1(new_n550), .B2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n592), .A2(new_n602), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  MUX2_X1   g181(.A(KEYINPUT81), .B(new_n604), .S(new_n606), .Z(G323));
  XOR2_X1   g182(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n608));
  XNOR2_X1  g183(.A(G323), .B(new_n608), .ZN(G282));
  NAND2_X1  g184(.A1(new_n472), .A2(new_n475), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n489), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n483), .A2(G123), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n619), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT83), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(KEYINPUT84), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(KEYINPUT84), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(G401));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT87), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(G229));
  MUX2_X1   g253(.A(G24), .B(G290), .S(G16), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1986), .ZN(new_n680));
  OR2_X1    g255(.A1(G25), .A2(G29), .ZN(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n682));
  INV_X1    g257(.A(G107), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G2105), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n483), .B2(G119), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n489), .A2(KEYINPUT89), .A3(G131), .ZN(new_n686));
  AOI21_X1  g261(.A(KEYINPUT89), .B1(new_n489), .B2(G131), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n681), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT35), .B(G1991), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n680), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT90), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n695), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G1971), .Z(new_n706));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n702), .A2(new_n703), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n694), .B1(new_n710), .B2(KEYINPUT34), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(KEYINPUT34), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n695), .A2(G19), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n550), .B2(new_n695), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT91), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1341), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  INV_X1    g294(.A(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G160), .B2(new_n689), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n695), .A2(G5), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G171), .B2(new_n695), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n689), .A2(G32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n489), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n732), .A2(new_n733), .B1(G105), .B2(new_n475), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n724), .B1(new_n726), .B2(G1961), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n718), .B1(KEYINPUT95), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n695), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n695), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT94), .B(G1966), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n689), .A2(G27), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT96), .Z(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n472), .A2(new_n497), .B1(new_n747), .B2(new_n495), .ZN(new_n748));
  INV_X1    g323(.A(new_n505), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n504), .B1(new_n472), .B2(new_n501), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n592), .B2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n755), .B1(new_n757), .B2(G1348), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n743), .B(new_n758), .C1(G1348), .C2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n695), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n489), .A2(G139), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  AOI22_X1  g341(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n766), .C1(new_n469), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n689), .A2(G33), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n772), .A2(G2072), .B1(G2084), .B2(new_n723), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT31), .B(G11), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G28), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n689), .B1(new_n775), .B2(G28), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .C1(new_n618), .C2(new_n689), .ZN(new_n778));
  INV_X1    g353(.A(G2072), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n771), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n736), .A2(new_n737), .B1(new_n726), .B2(G1961), .ZN(new_n781));
  AND4_X1   g356(.A1(new_n763), .A2(new_n773), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n739), .A2(new_n759), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n689), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n689), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n787), .B2(G2090), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G2090), .B2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n689), .A2(G26), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT28), .Z(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(G116), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G2105), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n483), .B2(G128), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n489), .A2(KEYINPUT92), .A3(G140), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT92), .B1(new_n489), .B2(G140), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n791), .B1(new_n802), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n783), .A2(new_n789), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n714), .A2(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  NAND2_X1  g383(.A1(new_n592), .A2(G559), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT38), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n518), .A2(G93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n512), .A2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n507), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n549), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n810), .B(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n817), .A2(new_n818), .A3(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(G145));
  AND2_X1   g397(.A1(new_n800), .A2(new_n801), .ZN(new_n823));
  NAND2_X1  g398(.A1(G164), .A2(KEYINPUT99), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n751), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n802), .A2(new_n827), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n489), .A2(G142), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n483), .A2(G130), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n834), .A2(new_n469), .A3(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n469), .B2(G118), .ZN(new_n836));
  OR2_X1    g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n835), .A2(G2104), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n831), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n829), .A2(new_n839), .A3(new_n830), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n688), .B(new_n611), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n768), .B(new_n735), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n491), .B(new_n618), .ZN(new_n850));
  XNOR2_X1  g425(.A(G160), .B(KEYINPUT98), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n848), .A2(KEYINPUT101), .A3(new_n849), .A4(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n848), .A2(new_n849), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(KEYINPUT102), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT40), .B1(new_n857), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(G395));
  XNOR2_X1  g438(.A(new_n815), .B(new_n605), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n565), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n592), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n565), .A2(new_n865), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n592), .A2(new_n865), .A3(new_n565), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n867), .A2(new_n868), .ZN(new_n875));
  INV_X1    g450(.A(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(KEYINPUT41), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n864), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT42), .ZN(new_n884));
  XOR2_X1   g459(.A(G290), .B(G305), .Z(new_n885));
  XOR2_X1   g460(.A(G303), .B(G288), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(KEYINPUT105), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n874), .B(new_n881), .C1(KEYINPUT105), .C2(new_n889), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n884), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n814), .A2(new_n594), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(G295));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n895), .ZN(G331));
  OR2_X1    g472(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(G168), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  NAND3_X1  g476(.A1(G171), .A2(new_n901), .A3(G286), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT106), .B1(G168), .B2(new_n539), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n815), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n815), .A2(new_n900), .A3(new_n902), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n879), .A3(new_n877), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n871), .A2(new_n906), .A3(new_n907), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n887), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT108), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n909), .A2(new_n913), .A3(new_n887), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n887), .B1(new_n909), .B2(new_n910), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n909), .A2(new_n910), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n887), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(KEYINPUT43), .A3(new_n916), .A4(new_n915), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g502(.A(G37), .B(new_n917), .C1(new_n912), .C2(new_n914), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n928), .B2(new_n920), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n919), .A2(new_n930), .A3(KEYINPUT43), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n920), .A3(new_n916), .A4(new_n915), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n927), .B1(new_n933), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n828), .B2(G1384), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n480), .A2(G2105), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n474), .A2(new_n937), .A3(G40), .A4(new_n476), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n823), .A2(new_n804), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n802), .A2(G2067), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n942), .B2(new_n735), .ZN(new_n943));
  NAND2_X1  g518(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n936), .A2(G1996), .A3(new_n938), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n939), .B(new_n946), .C1(KEYINPUT127), .C2(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n735), .B(new_n946), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n940), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n939), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n688), .B(new_n691), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n939), .ZN(new_n957));
  NOR2_X1   g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT110), .Z(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n939), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT48), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n954), .A2(new_n955), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n685), .B(new_n691), .C1(new_n686), .C2(new_n687), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n940), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n939), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NOR3_X1   g543(.A1(G164), .A2(new_n968), .A3(G1384), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n751), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n751), .A2(new_n970), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n938), .B1(KEYINPUT50), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1961), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(G164), .A2(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n938), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n754), .A2(KEYINPUT53), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n935), .A2(G1384), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n824), .A2(new_n826), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT114), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n824), .A2(new_n826), .A3(new_n986), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT113), .B(new_n935), .C1(G164), .C2(G1384), .ZN(new_n989));
  INV_X1    g564(.A(new_n938), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n975), .B2(new_n935), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n754), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n977), .B(new_n982), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n980), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n974), .A2(new_n1000), .A3(new_n976), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G286), .A2(G8), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(KEYINPUT51), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(KEYINPUT51), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n999), .B2(new_n1001), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1004), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1002), .A2(new_n1011), .B1(new_n1007), .B2(KEYINPUT51), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI211_X1 g589(.A(G301), .B(new_n997), .C1(new_n1014), .C2(KEYINPUT62), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n697), .A2(G1976), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n751), .A2(KEYINPUT115), .A3(new_n970), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n990), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(G8), .C1(G288), .C2(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1016), .A2(new_n1021), .A3(KEYINPUT52), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G305), .A2(G1981), .ZN(new_n1023));
  INV_X1    g598(.A(G1981), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n573), .A2(new_n574), .A3(new_n1024), .A4(new_n576), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(G8), .A3(new_n1019), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1022), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n994), .A2(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n974), .A2(new_n976), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G2090), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1035), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n973), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n938), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT50), .B1(new_n969), .B2(new_n971), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .A3(new_n990), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n978), .A2(new_n973), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n994), .A2(G1971), .B1(new_n1047), .B2(G2090), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1035), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT126), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1040), .A2(KEYINPUT126), .A3(new_n1049), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1015), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1010), .A2(G168), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1040), .A2(new_n1049), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(G8), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1034), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(KEYINPUT63), .A3(G168), .A4(new_n1010), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1055), .A2(KEYINPUT63), .B1(new_n1040), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1019), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1030), .A2(new_n1020), .A3(new_n697), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1009), .B(new_n1060), .C1(new_n1061), .C2(new_n1025), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1039), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(new_n1032), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1053), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1006), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n995), .A2(new_n996), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n477), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT125), .B1(new_n474), .B2(new_n476), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n937), .A2(KEYINPUT53), .A3(G40), .A4(new_n754), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n936), .A2(new_n988), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n977), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1068), .A2(G301), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n997), .B2(G301), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1066), .B1(new_n1067), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n997), .A2(G301), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1068), .A2(new_n1075), .A3(new_n1074), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(KEYINPUT54), .C1(new_n539), .C2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1078), .A2(new_n1050), .A3(new_n1051), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT118), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n565), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1047), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1047), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n994), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1088), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1088), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1083), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1037), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1060), .A2(new_n804), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n592), .ZN(new_n1106));
  INV_X1    g681(.A(new_n592), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1107), .A4(new_n1103), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1098), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1083), .B1(new_n1094), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1047), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1092), .B1(new_n1047), .B2(new_n1089), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1096), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1088), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1109), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n988), .A2(new_n946), .A3(new_n993), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1019), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT119), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1120), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1127), .B2(new_n550), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1120), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1119), .B(new_n550), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1118), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n550), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT120), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(KEYINPUT59), .A3(new_n1131), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1100), .A2(new_n1117), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1099), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1107), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1097), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1082), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n1140), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1065), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n939), .B1(new_n959), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT111), .Z(new_n1148));
  NAND4_X1  g723(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n967), .B1(new_n1145), .B2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g725(.A1(new_n639), .A2(new_n640), .ZN(new_n1152));
  NOR2_X1   g726(.A1(G227), .A2(new_n463), .ZN(new_n1153));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1153), .C1(new_n676), .C2(new_n677), .ZN(new_n1154));
  AOI21_X1  g728(.A(new_n1154), .B1(new_n857), .B2(new_n860), .ZN(new_n1155));
  AND2_X1   g729(.A1(new_n921), .A2(new_n926), .ZN(new_n1156));
  AND2_X1   g730(.A1(new_n1155), .A2(new_n1156), .ZN(G308));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(G225));
endmodule


