//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI211_X1 g035(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n464), .B2(G101), .ZN(new_n465));
  AND4_X1   g040(.A1(new_n462), .A2(new_n458), .A3(G101), .A4(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n459), .A2(new_n460), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n458), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G124), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G162));
  NAND2_X1  g056(.A1(KEYINPUT4), .A2(G138), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n458), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  AND2_X1   g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT69), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n498), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n502), .A2(new_n510), .ZN(G166));
  INV_X1    g086(.A(new_n504), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(G89), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n498), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n499), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n498), .A2(KEYINPUT70), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n524), .B2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT71), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n507), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(new_n534), .B2(new_n533), .ZN(new_n536));
  INV_X1    g111(.A(new_n509), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n524), .A2(G52), .B1(G90), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(new_n524), .A2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n507), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n509), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT74), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n499), .A2(KEYINPUT9), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n499), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n514), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n554), .A2(new_n555), .B1(G651), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n505), .A2(new_n498), .A3(G91), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(G299));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n537), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n500), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND3_X1  g144(.A1(new_n505), .A2(new_n498), .A3(G86), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n498), .A2(G48), .A3(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT77), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n512), .B2(new_n513), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n507), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n524), .A2(G47), .ZN(new_n579));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n514), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(G85), .A2(new_n537), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n524), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n522), .A2(KEYINPUT78), .A3(new_n523), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n587), .A2(G54), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n514), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT79), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n507), .B1(new_n592), .B2(KEYINPUT79), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n509), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n593), .A2(new_n594), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n585), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n585), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n562), .B(KEYINPUT76), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g188(.A(new_n472), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n464), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT80), .B(G2100), .Z(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n473), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n479), .A2(G123), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n619), .A2(new_n620), .A3(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n630), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  OR2_X1    g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT17), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  INV_X1    g225(.A(new_n647), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n645), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n650), .C1(new_n648), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n645), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT84), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  MUX2_X1   g252(.A(G19), .B(new_n545), .S(G16), .Z(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G1341), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n601), .A2(G16), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G4), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT87), .B(G1348), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n473), .A2(G140), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n479), .A2(G128), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n458), .A2(G116), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n686), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G29), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G26), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2067), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n679), .A2(new_n684), .A3(new_n685), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(G32), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n473), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G129), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n692), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT27), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1996), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n473), .A2(G139), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n614), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n458), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT89), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2072), .ZN(new_n721));
  NOR2_X1   g296(.A1(G27), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G164), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n709), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n692), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT24), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G34), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G160), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n730), .B1(new_n692), .B2(new_n625), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  INV_X1    g315(.A(G21), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G286), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G5), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G301), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n692), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n692), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n751), .B1(new_n754), .B2(G2090), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n726), .A2(new_n747), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT91), .B(KEYINPUT23), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT92), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n754), .A2(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n699), .B(new_n756), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G24), .ZN(new_n769));
  XNOR2_X1  g344(.A(G290), .B(KEYINPUT85), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1986), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n473), .A2(G131), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n479), .A2(G119), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n458), .A2(G107), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G25), .B(new_n777), .S(G29), .Z(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G23), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G288), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT33), .B(G1976), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G166), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G22), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g366(.A1(G6), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n577), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  INV_X1    g369(.A(G1981), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n781), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g374(.A(KEYINPUT86), .B(new_n798), .C1(new_n791), .C2(new_n796), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n791), .A2(new_n796), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(KEYINPUT34), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n799), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT36), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n799), .B(new_n806), .C1(new_n803), .C2(new_n800), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n768), .B1(new_n805), .B2(new_n807), .ZN(G311));
  XNOR2_X1  g383(.A(G311), .B(KEYINPUT94), .ZN(G150));
  AOI22_X1  g384(.A1(new_n524), .A2(G55), .B1(G93), .B2(new_n537), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(new_n507), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n546), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n812), .A2(new_n546), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n600), .A2(new_n608), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT96), .B(G860), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n812), .B2(new_n814), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n777), .B(KEYINPUT98), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(new_n616), .Z(new_n830));
  XOR2_X1   g405(.A(new_n496), .B(KEYINPUT97), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n716), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n705), .B(new_n690), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n479), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n458), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G142), .B2(new_n473), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n834), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n833), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n736), .B(new_n625), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G162), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(G37), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n842), .A2(KEYINPUT99), .A3(new_n845), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n841), .B2(new_n844), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g426(.A(G166), .B(G290), .ZN(new_n852));
  XNOR2_X1  g427(.A(G288), .B(new_n577), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT42), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(KEYINPUT103), .A3(new_n863), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n818), .B(new_n610), .ZN(new_n866));
  NAND2_X1  g441(.A1(G299), .A2(new_n601), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n605), .A2(new_n600), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n866), .B2(new_n869), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n864), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n864), .B1(new_n865), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(G868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n812), .A2(new_n814), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(G868), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G295));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n880), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  XNOR2_X1  g459(.A(G168), .B(G301), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n817), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(new_n815), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n818), .A2(new_n890), .A3(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n816), .A2(new_n817), .A3(new_n885), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n889), .A2(new_n891), .A3(new_n869), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n871), .B2(new_n872), .ZN(new_n895));
  INV_X1    g470(.A(new_n856), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n888), .A2(new_n869), .A3(new_n892), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(G299), .A2(new_n601), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n605), .A2(new_n600), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n870), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n869), .A2(new_n904), .A3(new_n870), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n889), .A2(new_n892), .A3(new_n891), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n884), .B(new_n897), .C1(new_n909), .C2(new_n896), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n883), .B1(new_n910), .B2(KEYINPUT43), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n907), .A2(new_n908), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n856), .B1(new_n912), .B2(new_n899), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n897), .A2(new_n884), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n915), .A3(KEYINPUT106), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n896), .B1(new_n893), .B2(new_n895), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n914), .A2(new_n918), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n910), .A2(new_n916), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n496), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n467), .ZN(new_n932));
  INV_X1    g507(.A(new_n470), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT107), .B(G40), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n705), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n690), .B(new_n696), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n779), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n777), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n690), .A2(G2067), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n937), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n777), .B(new_n779), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n937), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(G290), .A2(G1986), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT48), .B1(new_n936), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n936), .A2(KEYINPUT48), .A3(new_n949), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n936), .A2(new_n938), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT46), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT125), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(KEYINPUT46), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n940), .A2(new_n706), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n936), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n953), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  OR2_X1    g544(.A1(G288), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n496), .A2(G160), .A3(new_n928), .A4(new_n934), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(G8), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n970), .B(new_n971), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n929), .B2(new_n935), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(KEYINPUT113), .A3(new_n970), .A4(new_n971), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n970), .B1(new_n975), .B2(new_n976), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  OAI21_X1  g561(.A(G1981), .B1(new_n572), .B2(new_n576), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT77), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n573), .B(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G61), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n503), .B2(new_n504), .ZN(new_n992));
  OAI21_X1  g567(.A(G651), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(new_n795), .A3(new_n570), .A4(new_n571), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n987), .A2(new_n988), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT49), .B1(new_n995), .B2(KEYINPUT115), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n987), .A2(new_n994), .ZN(new_n997));
  NAND2_X1  g572(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n988), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n983), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n979), .A2(new_n984), .A3(new_n986), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT117), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n995), .A2(KEYINPUT115), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1000), .B1(new_n1005), .B2(KEYINPUT49), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n983), .A2(new_n1006), .B1(new_n985), .B2(KEYINPUT52), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n984), .A4(new_n979), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n1011));
  INV_X1    g586(.A(new_n935), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n931), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n931), .A2(KEYINPUT109), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n789), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n496), .A2(new_n1019), .A3(new_n928), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n496), .B2(new_n928), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n935), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1015), .A2(new_n1026), .A3(new_n789), .A4(new_n1016), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1018), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G303), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1031), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n935), .B1(new_n929), .B2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n1022), .B2(new_n935), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1021), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1024), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1017), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n974), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n738), .A3(new_n1020), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n496), .B2(new_n928), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n935), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1046), .B2(G1966), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n974), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G286), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1010), .A2(new_n1032), .A3(new_n1042), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1031), .B1(new_n1028), .B2(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1003), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1003), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1027), .A2(new_n1025), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1018), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT118), .B(new_n1056), .C1(new_n1059), .C2(new_n1031), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(KEYINPUT63), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1059), .B2(new_n1031), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1052), .A2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1006), .A2(G1976), .A3(G288), .ZN(new_n1065));
  INV_X1    g640(.A(new_n994), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n983), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1032), .B2(new_n1003), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1010), .A2(new_n1032), .A3(new_n1042), .ZN(new_n1069));
  AND2_X1   g644(.A1(G286), .A2(new_n974), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(KEYINPUT51), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1048), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1047), .A2(G286), .A3(new_n974), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT51), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1013), .A2(new_n744), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1057), .B1(new_n1075), .B2(new_n1043), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n1070), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT62), .B(new_n1072), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n724), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(G2078), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI221_X1 g659(.A(KEYINPUT123), .B1(new_n1013), .B2(new_n1084), .C1(new_n1023), .C2(G1961), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1013), .A2(new_n1084), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1961), .B1(new_n1034), .B2(new_n1020), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1078), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1073), .B(KEYINPUT51), .C1(new_n1070), .C2(new_n1076), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT62), .B1(new_n1093), .B2(new_n1072), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1068), .B1(new_n1069), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n562), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1097), .B(new_n1098), .C1(new_n559), .C2(new_n561), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1046), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1103), .B(new_n1105), .C1(new_n1038), .C2(G1956), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1038), .B2(G1956), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1103), .B(KEYINPUT121), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1034), .A2(new_n1020), .ZN(new_n1114));
  INV_X1    g689(.A(G1348), .ZN(new_n1115));
  INV_X1    g690(.A(new_n972), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1114), .A2(new_n1115), .B1(new_n696), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n600), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1107), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1103), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1108), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT61), .B1(new_n1122), .B2(new_n1106), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT122), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1117), .A2(new_n600), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT60), .B1(new_n1125), .B2(new_n1118), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT58), .B(G1341), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1013), .A2(G1996), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n546), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(new_n546), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1117), .A2(new_n1134), .A3(new_n601), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1106), .A2(KEYINPUT61), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1113), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1120), .B1(new_n1124), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1093), .A2(new_n1072), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1141));
  AND3_X1   g716(.A1(G160), .A2(G40), .A3(new_n1083), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1088), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1082), .A2(G301), .A3(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1081), .A2(new_n1080), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1140), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(G301), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1082), .A2(new_n1143), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1149), .B(KEYINPUT54), .C1(new_n1150), .C2(G301), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1069), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1064), .B(new_n1096), .C1(new_n1139), .C2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G290), .B(G1986), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n948), .B1(new_n936), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT108), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1153), .A2(KEYINPUT124), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n968), .B1(new_n1157), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g734(.A1(new_n659), .A2(G319), .ZN(new_n1161));
  NOR3_X1   g735(.A1(G229), .A2(G401), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g736(.A1(new_n920), .A2(new_n1162), .A3(new_n850), .ZN(G308));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n1162), .A3(new_n850), .ZN(G225));
endmodule


