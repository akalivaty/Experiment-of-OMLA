//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n483), .B1(new_n475), .B2(G136), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n463), .A2(new_n469), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(G164));
  AND2_X1   g072(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n499));
  OAI211_X1 g074(.A(KEYINPUT73), .B(G651), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n501), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(G651), .B1(new_n498), .B2(new_n499), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n515), .A2(new_n516), .B1(new_n504), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n510), .A2(G543), .A3(new_n500), .A4(new_n506), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT74), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n507), .A2(new_n510), .A3(new_n514), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  INV_X1    g099(.A(new_n521), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n517), .A2(new_n504), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT77), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n523), .B2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G51), .Z(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n519), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g114(.A(KEYINPUT76), .B(new_n535), .C1(new_n519), .C2(new_n536), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT78), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  AND2_X1   g120(.A1(new_n523), .A2(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n519), .A2(new_n547), .B1(new_n548), .B2(new_n504), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n515), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n519), .A2(new_n553), .B1(new_n554), .B2(new_n504), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT79), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n523), .A2(G91), .ZN(new_n563));
  INV_X1    g138(.A(new_n519), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .A3(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n519), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n504), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n563), .A2(new_n565), .A3(new_n568), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  AND2_X1   g148(.A1(new_n522), .A2(new_n528), .ZN(G303));
  NAND4_X1  g149(.A1(new_n507), .A2(G49), .A3(G543), .A4(new_n510), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n507), .A2(G87), .A3(new_n510), .A4(new_n514), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n513), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n523), .A2(G86), .B1(G651), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(G48), .A2(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n507), .A2(new_n510), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n507), .A2(KEYINPUT80), .A3(new_n510), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n582), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n589), .B1(new_n582), .B2(new_n588), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n519), .B2(new_n598), .C1(new_n515), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n504), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n519), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n515), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n605), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(G868), .B2(new_n610), .ZN(G284));
  OAI21_X1  g186(.A(new_n601), .B1(G868), .B2(new_n610), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G168), .B2(G868), .ZN(G280));
  XNOR2_X1  g189(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(new_n616), .B2(G860), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT83), .Z(G148));
  INV_X1    g193(.A(new_n610), .ZN(new_n619));
  OAI21_X1  g194(.A(G868), .B1(new_n619), .B2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g197(.A1(new_n463), .A2(new_n469), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(new_n473), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(KEYINPUT12), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(KEYINPUT12), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n475), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n460), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT84), .B(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT86), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n652), .B2(new_n655), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n664), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n664), .B(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n669), .B1(new_n671), .B2(new_n661), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n661), .A3(new_n665), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n667), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n689), .B(new_n688), .S(new_n681), .Z(new_n690));
  OR3_X1    g265(.A1(new_n687), .A2(new_n690), .A3(G1981), .ZN(new_n691));
  OAI21_X1  g266(.A(G1981), .B1(new_n687), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n692), .A3(G1986), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n695), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n678), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n677), .A3(new_n700), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(G34), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G160), .B2(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G2084), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G5), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G171), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n475), .A2(G141), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT97), .Z(new_n717));
  AND2_X1   g292(.A1(new_n473), .A2(G105), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT26), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n718), .B(new_n720), .C1(G129), .C2(new_n483), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(new_n707), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n707), .B2(G32), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n712), .B1(G1961), .B2(new_n715), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT100), .ZN(new_n728));
  NAND2_X1  g303(.A1(G299), .A2(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n713), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT23), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1956), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G139), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n476), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n623), .A2(G127), .ZN(new_n744));
  NAND2_X1  g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n460), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n743), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G29), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G33), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(G29), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2072), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n707), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n725), .B2(new_n726), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n707), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n483), .A2(G128), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(new_n707), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n707), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n707), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n711), .A2(G2084), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n758), .A2(new_n769), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n752), .A2(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n728), .A2(new_n734), .A3(new_n753), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n610), .B2(G16), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1348), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n713), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n556), .B2(new_n713), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1341), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n780), .A2(G1348), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n778), .A2(new_n781), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G286), .A2(new_n713), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1966), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1966), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT30), .B(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n707), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n635), .B2(new_n707), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n715), .B2(G1961), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n792), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n786), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G6), .B(G305), .S(G16), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n713), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n713), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(G1971), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(G1971), .ZN(new_n811));
  MUX2_X1   g386(.A(G23), .B(G288), .S(G16), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT33), .B(G1976), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n807), .A2(new_n818), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n707), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n483), .A2(G119), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT92), .Z(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G107), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n475), .B2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT93), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n822), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n831), .B2(new_n707), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n713), .A2(G24), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT94), .Z(new_n837));
  INV_X1    g412(.A(G290), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n713), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1986), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n817), .A2(new_n819), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n804), .B1(new_n843), .B2(new_n844), .ZN(G311));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n843), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(new_n802), .A3(new_n803), .A4(new_n786), .ZN(G150));
  INV_X1    g422(.A(new_n556), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n523), .A2(G93), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n564), .A2(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n513), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G651), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n849), .A2(new_n857), .A3(new_n850), .A4(new_n854), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n515), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n854), .B1(new_n519), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n856), .B1(new_n848), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n619), .A2(new_n616), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g444(.A(G860), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(G145));
  OAI21_X1  g449(.A(new_n722), .B1(new_n747), .B2(new_n749), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n746), .A2(new_n743), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n739), .B(KEYINPUT95), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n723), .A2(new_n876), .A3(new_n748), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n475), .A2(G142), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n483), .A2(G130), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n625), .A2(new_n626), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n627), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G164), .B(new_n765), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n831), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n828), .A2(new_n830), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n875), .A2(new_n878), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n888), .A2(new_n891), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n875), .B2(new_n878), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(new_n635), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G162), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n896), .A2(new_n900), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI211_X1 g484(.A(KEYINPUT102), .B(new_n902), .C1(new_n896), .C2(new_n900), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g487(.A(G303), .B1(new_n591), .B2(new_n592), .ZN(new_n913));
  XNOR2_X1  g488(.A(G290), .B(G288), .ZN(new_n914));
  INV_X1    g489(.A(new_n592), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(G166), .A3(new_n590), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n919), .A3(new_n916), .A4(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n916), .ZN(new_n922));
  INV_X1    g497(.A(new_n914), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT104), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  AOI211_X1 g500(.A(new_n925), .B(new_n914), .C1(new_n913), .C2(new_n916), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n864), .A2(new_n848), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n848), .A2(new_n855), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n619), .A2(G559), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n563), .A2(new_n568), .A3(new_n570), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n610), .A2(new_n565), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n610), .B1(new_n934), .B2(new_n565), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n619), .A2(G299), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n935), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n935), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n928), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n947), .A2(new_n928), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n864), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n952), .ZN(G295));
  OAI21_X1  g528(.A(new_n951), .B1(G868), .B2(new_n952), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n543), .A2(new_n544), .A3(G301), .ZN(new_n956));
  AOI21_X1  g531(.A(G301), .B1(new_n543), .B2(new_n544), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n956), .A2(new_n931), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G168), .A2(G171), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n543), .A2(new_n544), .A3(G301), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n865), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n942), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n931), .B1(new_n956), .B2(new_n957), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n865), .A3(new_n960), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n939), .A4(new_n935), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n922), .A2(new_n923), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n925), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n922), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n968), .A2(new_n969), .B1(new_n918), .B2(new_n920), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n904), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n944), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n942), .B2(KEYINPUT106), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n958), .A2(new_n961), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n955), .B(new_n971), .C1(new_n970), .C2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n966), .A2(new_n970), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT44), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n971), .B2(new_n977), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n970), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n927), .A2(new_n962), .A3(new_n965), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n955), .A3(new_n983), .A4(new_n904), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n980), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(new_n478), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n470), .A2(new_n471), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n989), .B(G40), .C1(new_n990), .C2(new_n460), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n722), .B(G1996), .Z(new_n995));
  XNOR2_X1  g570(.A(new_n765), .B(new_n768), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n892), .A2(new_n834), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n892), .A2(new_n834), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(G290), .B(G1986), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT62), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  INV_X1    g580(.A(G1966), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n472), .A2(new_n478), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(new_n993), .A3(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n494), .A2(new_n496), .ZN(new_n1010));
  INV_X1    g585(.A(new_n491), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT116), .B1(new_n1008), .B2(new_n993), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT117), .B(new_n1006), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT108), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2084), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n991), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1021), .A2(new_n1024), .A3(new_n1027), .A4(new_n1022), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1016), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1008), .A2(new_n993), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n1013), .A3(new_n1009), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1006), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1029), .A2(G286), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1005), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1033), .A2(new_n1006), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(G168), .A3(new_n1041), .A4(new_n1016), .ZN(new_n1042));
  OAI21_X1  g617(.A(G286), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1037), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1004), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1037), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(KEYINPUT62), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(KEYINPUT109), .A3(G8), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n582), .A2(new_n588), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n582), .B2(new_n588), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n582), .A2(new_n588), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G1981), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n1060), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1058), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT113), .B(new_n1058), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n575), .A2(new_n576), .A3(G1976), .A4(new_n577), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1058), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1056), .A2(new_n1057), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1085), .B(KEYINPUT112), .Z(new_n1086));
  AOI22_X1  g661(.A1(new_n1079), .A2(new_n1083), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n522), .A2(new_n528), .A3(G8), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT55), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1008), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1092), .A2(KEYINPUT115), .ZN(new_n1093));
  AOI21_X1  g668(.A(G2090), .B1(new_n1092), .B2(KEYINPUT115), .ZN(new_n1094));
  INV_X1    g669(.A(G1971), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1013), .A2(new_n1008), .A3(new_n993), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1093), .A2(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1089), .B1(new_n1036), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(new_n1088), .B(KEYINPUT55), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1095), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT107), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(KEYINPUT107), .A3(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(G2090), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(G8), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1072), .A2(new_n1087), .A3(new_n1098), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1961), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n772), .A2(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1096), .B2(G2078), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI221_X1 g690(.A(new_n1109), .B1(new_n1033), .B2(new_n1110), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1107), .A2(G301), .A3(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1048), .A2(new_n1052), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1105), .A2(G8), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n1089), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1072), .A2(new_n1087), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1060), .B(KEYINPUT114), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G288), .A2(G1976), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1072), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1058), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1122), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G286), .A2(new_n1036), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1107), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1129), .B(KEYINPUT63), .C1(new_n1029), .C2(new_n1034), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1120), .A2(KEYINPUT119), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1099), .B1(new_n1120), .B2(KEYINPUT119), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(new_n1106), .A3(new_n1072), .A4(new_n1087), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1053), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(G1996), .B2(new_n1096), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT59), .A4(new_n556), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n556), .B1(new_n1138), .B2(KEYINPUT59), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1092), .A2(new_n733), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT56), .B(G2072), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1096), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  NAND3_X1  g724(.A1(G299), .A2(new_n1149), .A3(KEYINPUT57), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(G299), .B2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(G299), .A2(new_n1149), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1096), .A2(new_n1147), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1150), .A4(new_n1145), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1158), .A3(KEYINPUT61), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1144), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1156), .A2(new_n1150), .B1(new_n1157), .B2(new_n1145), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1053), .A2(G2067), .ZN(new_n1167));
  INV_X1    g742(.A(G1348), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1104), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n619), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n619), .B1(new_n1169), .B2(KEYINPUT60), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1170), .A2(new_n1171), .B1(KEYINPUT60), .B2(new_n1169), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT123), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1160), .A2(new_n1166), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1153), .B1(new_n1169), .B2(new_n619), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1158), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G171), .B(KEYINPUT54), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1109), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1096), .B2(new_n1110), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1117), .A2(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1107), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1179), .A2(new_n1184), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1137), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1003), .B1(new_n1119), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n994), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n998), .B1(new_n997), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(G2067), .B2(new_n765), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1190), .A2(KEYINPUT126), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(KEYINPUT126), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n994), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1188), .B1(new_n996), .B2(new_n723), .ZN(new_n1194));
  OR3_X1    g769(.A1(new_n1188), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT46), .B1(new_n1188), .B2(G1996), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT47), .Z(new_n1198));
  NAND2_X1  g773(.A1(new_n1001), .A2(new_n994), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n838), .A2(new_n994), .A3(new_n694), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1201), .A2(KEYINPUT48), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(KEYINPUT48), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1193), .A2(new_n1198), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1187), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n658), .A2(G319), .ZN(new_n1209));
  OR2_X1    g783(.A1(new_n1209), .A2(G227), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n703), .B2(new_n705), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n911), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1208), .B1(new_n985), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g788(.A(KEYINPUT127), .B(new_n1212), .C1(new_n981), .C2(new_n984), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1214), .A2(new_n1215), .ZN(G308));
  NAND2_X1  g790(.A1(new_n985), .A2(new_n1213), .ZN(G225));
endmodule


