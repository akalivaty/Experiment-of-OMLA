

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n724), .ZN(n705) );
  BUF_X1 U549 ( .A(n612), .Z(n613) );
  BUF_X1 U550 ( .A(n608), .Z(n609) );
  AND2_X2 U551 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NOR2_X1 U552 ( .A1(n805), .A2(n804), .ZN(n514) );
  XOR2_X1 U553 ( .A(KEYINPUT32), .B(KEYINPUT100), .Z(n515) );
  XOR2_X1 U554 ( .A(G543), .B(KEYINPUT0), .Z(n516) );
  OR2_X1 U555 ( .A1(n771), .A2(n770), .ZN(n517) );
  XNOR2_X1 U556 ( .A(n766), .B(KEYINPUT105), .ZN(n518) );
  OR2_X1 U557 ( .A1(n918), .A2(n701), .ZN(n702) );
  NOR2_X1 U558 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U559 ( .A1(n773), .A2(n681), .ZN(n724) );
  NAND2_X1 U560 ( .A1(G160), .A2(G40), .ZN(n772) );
  INV_X1 U561 ( .A(KEYINPUT13), .ZN(n566) );
  NOR2_X1 U562 ( .A1(n549), .A2(n653), .ZN(n647) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n646) );
  XNOR2_X1 U564 ( .A(n567), .B(n566), .ZN(n568) );
  NOR2_X1 U565 ( .A1(G651), .A2(n653), .ZN(n658) );
  NAND2_X1 U566 ( .A1(n571), .A2(n570), .ZN(n927) );
  NOR2_X1 U567 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U568 ( .A1(G113), .A2(n894), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n519), .B(KEYINPUT64), .ZN(n522) );
  INV_X1 U570 ( .A(G2104), .ZN(n525) );
  NOR2_X2 U571 ( .A1(G2105), .A2(n525), .ZN(n608) );
  NAND2_X1 U572 ( .A1(G101), .A2(n608), .ZN(n520) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U574 ( .A1(n522), .A2(n521), .ZN(n529) );
  XNOR2_X1 U575 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U577 ( .A(n524), .B(n523), .ZN(n612) );
  NAND2_X1 U578 ( .A1(G137), .A2(n612), .ZN(n527) );
  AND2_X1 U579 ( .A1(n525), .A2(G2105), .ZN(n893) );
  NAND2_X1 U580 ( .A1(G125), .A2(n893), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U582 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U583 ( .A(G82), .ZN(G220) );
  INV_X1 U584 ( .A(G132), .ZN(G219) );
  INV_X1 U585 ( .A(G108), .ZN(G238) );
  INV_X1 U586 ( .A(G69), .ZN(G235) );
  INV_X1 U587 ( .A(G120), .ZN(G236) );
  NOR2_X1 U588 ( .A1(G220), .A2(G219), .ZN(n530) );
  XOR2_X1 U589 ( .A(KEYINPUT22), .B(n530), .Z(n531) );
  NOR2_X1 U590 ( .A1(G218), .A2(n531), .ZN(n532) );
  XNOR2_X1 U591 ( .A(KEYINPUT82), .B(n532), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n533), .A2(G96), .ZN(n840) );
  NAND2_X1 U593 ( .A1(n840), .A2(G2106), .ZN(n538) );
  NOR2_X1 U594 ( .A1(G235), .A2(G236), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n534), .B(KEYINPUT83), .ZN(n535) );
  NOR2_X1 U596 ( .A1(G238), .A2(n535), .ZN(n536) );
  NAND2_X1 U597 ( .A1(G57), .A2(n536), .ZN(n841) );
  NAND2_X1 U598 ( .A1(n841), .A2(G567), .ZN(n537) );
  AND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(G319) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(G138), .A2(n612), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G102), .A2(n608), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G126), .A2(n893), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G114), .A2(n894), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(G164) );
  NAND2_X1 U608 ( .A1(n646), .A2(G89), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT4), .ZN(n547) );
  INV_X1 U610 ( .A(G651), .ZN(n549) );
  XNOR2_X1 U611 ( .A(KEYINPUT66), .B(n516), .ZN(n653) );
  NAND2_X1 U612 ( .A1(G76), .A2(n647), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT5), .ZN(n555) );
  NOR2_X1 U615 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U616 ( .A(KEYINPUT1), .B(n550), .Z(n657) );
  NAND2_X1 U617 ( .A1(G63), .A2(n657), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G51), .A2(n658), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U624 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n558) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n836) );
  NAND2_X1 U628 ( .A1(n836), .A2(G567), .ZN(n559) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U630 ( .A1(G56), .A2(n657), .ZN(n560) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n560), .Z(n569) );
  NAND2_X1 U632 ( .A1(n647), .A2(G68), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n562) );
  NAND2_X1 U634 ( .A1(G81), .A2(n646), .ZN(n561) );
  XNOR2_X1 U635 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U636 ( .A(KEYINPUT72), .B(n563), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n567) );
  NOR2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n658), .A2(G43), .ZN(n570) );
  INV_X1 U640 ( .A(G860), .ZN(n601) );
  OR2_X1 U641 ( .A1(n927), .A2(n601), .ZN(G153) );
  XNOR2_X1 U642 ( .A(KEYINPUT9), .B(KEYINPUT69), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G90), .A2(n646), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G77), .A2(n647), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U646 ( .A(n575), .B(n574), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n657), .A2(G64), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT68), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G52), .A2(n658), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G171) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G301), .A2(G868), .ZN(n581) );
  XNOR2_X1 U654 ( .A(n581), .B(KEYINPUT74), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G66), .A2(n657), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G92), .A2(n646), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G54), .A2(n658), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G79), .A2(n647), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U662 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n588) );
  XNOR2_X1 U663 ( .A(n589), .B(n588), .ZN(n918) );
  OR2_X1 U664 ( .A1(G868), .A2(n918), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G65), .A2(n657), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G78), .A2(n647), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n646), .A2(G91), .ZN(n594) );
  XOR2_X1 U670 ( .A(KEYINPUT70), .B(n594), .Z(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n658), .A2(G53), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(G299) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n600) );
  INV_X1 U675 ( .A(G868), .ZN(n671) );
  NOR2_X1 U676 ( .A1(G286), .A2(n671), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n602), .A2(n918), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n927), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G868), .A2(n918), .ZN(n604) );
  NOR2_X1 U683 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G282) );
  XOR2_X1 U685 ( .A(G2100), .B(KEYINPUT76), .Z(n619) );
  NAND2_X1 U686 ( .A1(G123), .A2(n893), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n609), .A2(G99), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G135), .A2(n613), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G111), .A2(n894), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n991) );
  XNOR2_X1 U694 ( .A(G2096), .B(n991), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n918), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(n927), .ZN(n668) );
  NOR2_X1 U698 ( .A1(n668), .A2(G860), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G67), .A2(n657), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G93), .A2(n646), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G55), .A2(n658), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G80), .A2(n647), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n670) );
  XOR2_X1 U706 ( .A(n627), .B(n670), .Z(G145) );
  NAND2_X1 U707 ( .A1(G61), .A2(n657), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G86), .A2(n646), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n647), .A2(G73), .ZN(n630) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n658), .A2(G48), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G88), .A2(n646), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G62), .A2(n657), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G50), .A2(n658), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G75), .A2(n647), .ZN(n637) );
  XNOR2_X1 U720 ( .A(KEYINPUT79), .B(n637), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT80), .ZN(G303) );
  NAND2_X1 U724 ( .A1(n658), .A2(G47), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n657), .A2(G60), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U727 ( .A(KEYINPUT67), .B(n645), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G85), .A2(n646), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G72), .A2(n647), .ZN(n648) );
  AND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(G290) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(KEYINPUT78), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G87), .A2(n653), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G49), .A2(n658), .ZN(n659) );
  XOR2_X1 U738 ( .A(KEYINPUT77), .B(n659), .Z(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(G288) );
  XNOR2_X1 U740 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n663) );
  INV_X1 U741 ( .A(G299), .ZN(n915) );
  XNOR2_X1 U742 ( .A(G305), .B(n915), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n665) );
  XNOR2_X1 U744 ( .A(G303), .B(G290), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n665), .B(n664), .ZN(n667) );
  XOR2_X1 U746 ( .A(G288), .B(n670), .Z(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n905) );
  XNOR2_X1 U748 ( .A(n668), .B(n905), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n677), .A2(G2072), .ZN(G158) );
  NAND2_X1 U757 ( .A1(G661), .A2(G483), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT84), .B(n678), .Z(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G319), .ZN(n680) );
  XNOR2_X1 U760 ( .A(n680), .B(KEYINPUT85), .ZN(n839) );
  NAND2_X1 U761 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U763 ( .A(KEYINPUT94), .B(G1961), .ZN(n941) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n773) );
  INV_X1 U765 ( .A(n772), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n941), .A2(n724), .ZN(n683) );
  XOR2_X1 U767 ( .A(G2078), .B(KEYINPUT25), .Z(n973) );
  NAND2_X1 U768 ( .A1(n705), .A2(n973), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U770 ( .A(n684), .B(KEYINPUT95), .Z(n716) );
  AND2_X1 U771 ( .A1(G301), .A2(n716), .ZN(n689) );
  NAND2_X1 U772 ( .A1(G8), .A2(n724), .ZN(n771) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n771), .ZN(n738) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n724), .ZN(n734) );
  NOR2_X1 U775 ( .A1(n738), .A2(n734), .ZN(n685) );
  NAND2_X1 U776 ( .A1(G8), .A2(n685), .ZN(n686) );
  XNOR2_X1 U777 ( .A(KEYINPUT30), .B(n686), .ZN(n687) );
  NOR2_X1 U778 ( .A1(G168), .A2(n687), .ZN(n688) );
  NOR2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U780 ( .A(KEYINPUT31), .B(n690), .ZN(n720) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n705), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT26), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G1341), .A2(n724), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n695) );
  INV_X1 U785 ( .A(KEYINPUT97), .ZN(n694) );
  XNOR2_X1 U786 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n696), .A2(n927), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n701), .A2(n918), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n705), .A2(G1348), .ZN(n698) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n724), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n709) );
  NAND2_X1 U794 ( .A1(n705), .A2(G2072), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n704), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U796 ( .A(G1956), .ZN(n942) );
  NOR2_X1 U797 ( .A1(n942), .A2(n705), .ZN(n706) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n710), .A2(n915), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U801 ( .A1(n710), .A2(n915), .ZN(n712) );
  XOR2_X1 U802 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n711) );
  XNOR2_X1 U803 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n715), .B(KEYINPUT29), .ZN(n718) );
  NOR2_X1 U806 ( .A1(G301), .A2(n716), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n719) );
  INV_X1 U808 ( .A(KEYINPUT98), .ZN(n721) );
  XNOR2_X1 U809 ( .A(n722), .B(n721), .ZN(n736) );
  AND2_X1 U810 ( .A1(G286), .A2(G8), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n736), .A2(n723), .ZN(n732) );
  INV_X1 U812 ( .A(G8), .ZN(n730) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n771), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U816 ( .A1(G303), .A2(n727), .ZN(n728) );
  XOR2_X1 U817 ( .A(KEYINPUT99), .B(n728), .Z(n729) );
  OR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U820 ( .A(n733), .B(n515), .ZN(n742) );
  NAND2_X1 U821 ( .A1(G8), .A2(n734), .ZN(n735) );
  XOR2_X1 U822 ( .A(KEYINPUT93), .B(n735), .Z(n740) );
  INV_X1 U823 ( .A(n736), .ZN(n737) );
  NOR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n751) );
  NAND2_X1 U827 ( .A1(G8), .A2(G166), .ZN(n743) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n743), .ZN(n744) );
  XNOR2_X1 U829 ( .A(n744), .B(KEYINPUT103), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n751), .A2(n745), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT104), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n747), .A2(n771), .ZN(n765) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U834 ( .A1(G303), .A2(G1971), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n755), .A2(n748), .ZN(n934) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n749) );
  AND2_X1 U837 ( .A1(n934), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n762) );
  INV_X1 U839 ( .A(n771), .ZN(n753) );
  NAND2_X1 U840 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XOR2_X1 U841 ( .A(KEYINPUT101), .B(n752), .Z(n921) );
  AND2_X1 U842 ( .A1(n753), .A2(n921), .ZN(n754) );
  OR2_X1 U843 ( .A1(KEYINPUT33), .A2(n754), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n756), .A2(n771), .ZN(n758) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n923) );
  INV_X1 U847 ( .A(n923), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(n763), .B(KEYINPUT102), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U853 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n767) );
  XNOR2_X1 U854 ( .A(n767), .B(KEYINPUT91), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XNOR2_X1 U856 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n518), .A2(n517), .ZN(n806) );
  NOR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n820) );
  NAND2_X1 U859 ( .A1(G140), .A2(n613), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G104), .A2(n609), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n776), .ZN(n783) );
  NAND2_X1 U863 ( .A1(n893), .A2(G128), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT86), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G116), .A2(n894), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT87), .B(n780), .ZN(n781) );
  XNOR2_X1 U868 ( .A(KEYINPUT35), .B(n781), .ZN(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT36), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT88), .ZN(n880) );
  XNOR2_X1 U872 ( .A(KEYINPUT37), .B(G2067), .ZN(n818) );
  NOR2_X1 U873 ( .A1(n880), .A2(n818), .ZN(n998) );
  NAND2_X1 U874 ( .A1(n820), .A2(n998), .ZN(n817) );
  INV_X1 U875 ( .A(n817), .ZN(n805) );
  NAND2_X1 U876 ( .A1(G141), .A2(n613), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G129), .A2(n893), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n609), .A2(G105), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n894), .A2(G117), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n878) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n878), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G95), .A2(n609), .ZN(n793) );
  XNOR2_X1 U886 ( .A(n793), .B(KEYINPUT90), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G131), .A2(n613), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G119), .A2(n893), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G107), .A2(n894), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT89), .B(n796), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n877) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n877), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n994) );
  NAND2_X1 U896 ( .A1(n820), .A2(n994), .ZN(n808) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n936) );
  NAND2_X1 U898 ( .A1(n820), .A2(n936), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n808), .A2(n803), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n806), .A2(n514), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(KEYINPUT106), .ZN(n823) );
  XOR2_X1 U902 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n815) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n878), .ZN(n989) );
  INV_X1 U904 ( .A(n808), .ZN(n811) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n877), .ZN(n992) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n992), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n989), .A2(n812), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT107), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n880), .A2(n818), .ZN(n1009) );
  NAND2_X1 U914 ( .A1(n819), .A2(n1009), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U918 ( .A(G2435), .B(G2443), .ZN(n834) );
  XOR2_X1 U919 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n826) );
  XNOR2_X1 U920 ( .A(G2454), .B(G2430), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U922 ( .A(G2427), .B(G2438), .Z(n828) );
  XNOR2_X1 U923 ( .A(G1348), .B(G1341), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U925 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U926 ( .A(G2446), .B(G2451), .ZN(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(G14), .ZN(n909) );
  XNOR2_X1 U930 ( .A(KEYINPUT111), .B(n909), .ZN(G401) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(G1956), .B(KEYINPUT41), .ZN(n851) );
  XOR2_X1 U941 ( .A(G1971), .B(G1966), .Z(n843) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1961), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(G1976), .B(G1986), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT112), .B(G2474), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U951 ( .A(G2096), .B(G2100), .Z(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2090), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U960 ( .A1(G124), .A2(n893), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n609), .A2(G100), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G136), .A2(n613), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G112), .A2(n894), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U968 ( .A1(n894), .A2(G118), .ZN(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT113), .B(n867), .ZN(n876) );
  XOR2_X1 U970 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT45), .B(n868), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G142), .A2(n613), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G106), .A2(n609), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G130), .A2(n893), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n882) );
  XOR2_X1 U979 ( .A(n878), .B(n877), .Z(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n885) );
  XNOR2_X1 U982 ( .A(G164), .B(G162), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n883), .B(n991), .ZN(n884) );
  XOR2_X1 U984 ( .A(n885), .B(n884), .Z(n890) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(n888), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n901) );
  NAND2_X1 U990 ( .A1(G139), .A2(n613), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G103), .A2(n609), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G127), .A2(n893), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n1002) );
  XNOR2_X1 U998 ( .A(n1002), .B(G160), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n927), .B(KEYINPUT119), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(G171), .B(n918), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n905), .B(G286), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(G397) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .ZN(n940) );
  XNOR2_X1 U1016 ( .A(n915), .B(G1956), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1019 ( .A(G1348), .B(n918), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G168), .B(G1966), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT124), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT57), .B(n926), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(G301), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n927), .B(G1341), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n938) );
  INV_X1 U1031 ( .A(n934), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n1018) );
  XOR2_X1 U1035 ( .A(n941), .B(G5), .Z(n952) );
  XNOR2_X1 U1036 ( .A(G20), .B(n942), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G19), .B(G1341), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT59), .B(G1348), .Z(n947) );
  XNOR2_X1 U1042 ( .A(G4), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n950), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n963) );
  XOR2_X1 U1046 ( .A(G1966), .B(G21), .Z(n961) );
  XOR2_X1 U1047 ( .A(G1971), .B(G22), .Z(n955) );
  XOR2_X1 U1048 ( .A(G24), .B(KEYINPUT126), .Z(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(G1986), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT125), .B(G1976), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G23), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT58), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G11), .ZN(n1016) );
  XOR2_X1 U1061 ( .A(G34), .B(KEYINPUT122), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G2084), .B(KEYINPUT54), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n984) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n982) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G26), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G32), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G27), .B(n973), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(G29), .A2(n986), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT55), .ZN(n1014) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1083 ( .A(KEYINPUT51), .B(n990), .Z(n1000) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n996) );
  XOR2_X1 U1085 ( .A(G160), .B(G2084), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT120), .B(n1001), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G2072), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G164), .B(G2078), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT121), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(G29), .A2(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

