//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n207), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n214), .B(new_n217), .C1(new_n220), .C2(new_n223), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n202), .A2(G68), .ZN(new_n238));
  INV_X1    g0038(.A(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n237), .B(new_n243), .ZN(G351));
  AOI21_X1  g0044(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT71), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT71), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n251), .C2(new_n246), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G238), .ZN(new_n256));
  OR3_X1    g0056(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G226), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G232), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(G1698), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G97), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n251), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n245), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n245), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n248), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n257), .A2(new_n268), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n261), .A2(new_n264), .B1(G33), .B2(G97), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(new_n252), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT13), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n257), .A2(new_n268), .A3(new_n272), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G169), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n273), .A2(new_n277), .A3(G179), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n279), .A2(new_n281), .A3(new_n285), .A4(G169), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n239), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n251), .A2(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n218), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT12), .B1(new_n300), .B2(G68), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT12), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n239), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n239), .B1(new_n253), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n298), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .A4(new_n307), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n287), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n280), .B2(KEYINPUT13), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n273), .B1(new_n310), .B2(new_n311), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n279), .A2(G200), .A3(new_n281), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT74), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n258), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G33), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(G226), .A2(G1698), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n260), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT78), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT78), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(new_n328), .A3(new_n260), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n324), .A2(G223), .A3(new_n331), .A4(new_n260), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n327), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n245), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n252), .A2(new_n254), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n252), .A2(G274), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n263), .A2(new_n335), .B1(new_n336), .B2(new_n254), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(G179), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n333), .B2(new_n245), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n251), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT7), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(G20), .ZN(new_n349));
  AOI21_X1  g0149(.A(G33), .B1(new_n322), .B2(new_n323), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n347), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n261), .B2(G20), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n239), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G58), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n239), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(new_n201), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n343), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(G20), .B1(new_n324), .B2(new_n260), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n361), .B2(new_n348), .ZN(new_n362));
  AOI211_X1 g0162(.A(KEYINPUT7), .B(G20), .C1(new_n324), .C2(new_n260), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT16), .B(new_n358), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n295), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n300), .ZN(new_n367));
  INV_X1    g0167(.A(new_n295), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n300), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT67), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT67), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n305), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n370), .A2(new_n372), .B1(new_n253), .B2(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n373), .B2(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n342), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT18), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n334), .B2(new_n338), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n314), .B(new_n337), .C1(new_n333), .C2(new_n245), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n365), .A4(new_n374), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n342), .A2(new_n375), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n334), .A2(G190), .A3(new_n338), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n378), .B2(new_n341), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n387), .B2(new_n375), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n377), .A2(new_n382), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT79), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G222), .A2(G1698), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n331), .A2(G223), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n261), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n245), .C1(G77), .C2(new_n261), .ZN(new_n395));
  INV_X1    g0195(.A(new_n335), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G226), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(new_n272), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n314), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(G200), .B2(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n300), .A2(new_n202), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n373), .B2(new_n202), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT68), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT68), .B(new_n402), .C1(new_n373), .C2(new_n202), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n366), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n290), .B1(G150), .B2(new_n288), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n203), .A2(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n368), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n401), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(KEYINPUT9), .B(new_n411), .C1(new_n405), .C2(new_n406), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n400), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT10), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT10), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n400), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n398), .A2(G179), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n407), .A2(new_n412), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n398), .A2(new_n340), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(G77), .B1(new_n219), .B2(G1), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n369), .A2(new_n426), .B1(G77), .B2(new_n300), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n408), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT15), .B(G87), .Z(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n291), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n431), .B2(new_n295), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G244), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n272), .B1(new_n434), .B2(new_n335), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n261), .A2(G232), .A3(new_n331), .ZN(new_n437));
  INV_X1    g0237(.A(G107), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n261), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n435), .B1(new_n439), .B2(new_n245), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(G169), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(KEYINPUT70), .B(new_n432), .C1(new_n440), .C2(new_n378), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(G190), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n432), .B1(new_n440), .B2(new_n378), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT70), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n419), .A2(new_n425), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n390), .A2(KEYINPUT79), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n320), .A2(new_n391), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n239), .A2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n324), .A2(new_n260), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n291), .B2(new_n266), .ZN(new_n459));
  NAND3_X1  g0259(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n219), .ZN(new_n461));
  INV_X1    g0261(.A(G87), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n266), .A3(new_n438), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT83), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n457), .B(new_n459), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n463), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n457), .A4(new_n459), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(new_n474), .A3(new_n295), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n430), .A2(new_n302), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n253), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n368), .A2(new_n300), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n478), .A2(new_n480), .B1(G87), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT82), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n247), .A2(G1), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(new_n252), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n485), .A3(new_n252), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(new_n271), .B2(new_n486), .ZN(new_n492));
  INV_X1    g0292(.A(new_n260), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n345), .A2(new_n346), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G33), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G238), .A2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n434), .B2(G1698), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n495), .A2(new_n497), .B1(G33), .B2(G116), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n492), .B(new_n314), .C1(new_n252), .C2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n252), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n271), .A2(new_n486), .ZN(new_n501));
  INV_X1    g0301(.A(new_n491), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n489), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n499), .B1(new_n504), .B2(G200), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n482), .A2(new_n430), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n479), .B1(new_n475), .B2(new_n476), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n442), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n340), .B1(new_n500), .B2(new_n503), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n484), .A2(new_n505), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n294), .A2(new_n218), .B1(G20), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n219), .C1(G33), .C2(new_n266), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(KEYINPUT20), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT20), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n302), .A2(new_n516), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n482), .B2(new_n516), .ZN(new_n524));
  OAI21_X1  g0324(.A(G169), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT5), .B(G41), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(new_n252), .A3(G274), .A4(new_n486), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n486), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n252), .ZN(new_n529));
  INV_X1    g0329(.A(G270), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G257), .A2(G1698), .ZN(new_n532));
  INV_X1    g0332(.A(G264), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(G1698), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n324), .A3(new_n260), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n259), .A2(new_n260), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G303), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n252), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n515), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n245), .B1(new_n486), .B2(new_n526), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G270), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n495), .A2(new_n534), .B1(G303), .B2(new_n536), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n527), .B(new_n542), .C1(new_n543), .C2(new_n252), .ZN(new_n544));
  OAI221_X1 g0344(.A(new_n523), .B1(new_n482), .B2(new_n516), .C1(new_n520), .C2(new_n521), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT21), .A4(G169), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(new_n545), .A3(G179), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n544), .B2(G200), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n314), .B2(new_n544), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n462), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n324), .A2(new_n260), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n219), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n219), .A2(G87), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n555), .B1(new_n536), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT23), .B1(new_n219), .B2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT86), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n219), .C2(G107), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n219), .A2(KEYINPUT23), .A3(G107), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n562), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n554), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(new_n557), .B2(new_n558), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n562), .A2(new_n567), .A3(new_n568), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT24), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n295), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT25), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n300), .B2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n300), .A2(new_n575), .A3(G107), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n482), .A2(new_n438), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  MUX2_X1   g0381(.A(G250), .B(G257), .S(G1698), .Z(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n324), .A3(new_n260), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n252), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n541), .A2(G264), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n527), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n442), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(G200), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n585), .B1(G264), .B2(new_n541), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(G190), .A3(new_n527), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n574), .A2(new_n592), .A3(new_n580), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n438), .B1(new_n352), .B2(new_n353), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n288), .A2(G77), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n599), .A2(new_n266), .A3(G107), .ZN(new_n600));
  XNOR2_X1  g0400(.A(G97), .B(G107), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n602), .B2(new_n219), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n295), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT80), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n300), .B2(G97), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n302), .A2(KEYINPUT80), .A3(new_n266), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n483), .A2(G97), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n324), .A2(new_n260), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n434), .A2(G1698), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n259), .A2(new_n260), .A3(G250), .A4(G1698), .ZN(new_n615));
  AND2_X1   g0415(.A1(KEYINPUT4), .A2(G244), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n259), .A2(new_n260), .A3(new_n616), .A4(new_n331), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n615), .A2(new_n617), .A3(new_n518), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n252), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n528), .A2(G257), .A3(new_n252), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n527), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n340), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT4), .B1(new_n495), .B2(new_n612), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n615), .A2(new_n617), .A3(new_n518), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n245), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n621), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n442), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n609), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n619), .B2(new_n621), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT81), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n614), .A2(new_n618), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n621), .B1(new_n631), .B2(new_n245), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n629), .A2(new_n630), .B1(new_n632), .B2(G190), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n625), .A2(new_n630), .A3(G190), .A4(new_n626), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n604), .A3(new_n608), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n628), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n596), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n455), .A2(new_n514), .A3(new_n553), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n512), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(KEYINPUT87), .B(new_n340), .C1(new_n500), .C2(new_n503), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n640), .A2(new_n511), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n510), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n595), .B(new_n628), .C1(new_n633), .C2(new_n635), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n548), .B1(new_n590), .B2(new_n581), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n483), .A2(G87), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n648), .B(new_n505), .C1(new_n508), .C2(new_n509), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n628), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n506), .B1(new_n478), .B2(new_n480), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n640), .A2(new_n511), .A3(new_n641), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n649), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n510), .A2(new_n513), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n649), .A4(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n454), .B1(new_n650), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n444), .ZN(new_n661));
  INV_X1    g0461(.A(new_n318), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n313), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n382), .A2(new_n388), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n342), .A2(new_n375), .A3(new_n383), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n383), .B1(new_n342), .B2(new_n375), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n419), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n425), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n660), .A2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n253), .A2(new_n219), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n545), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n552), .B2(KEYINPUT88), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(KEYINPUT88), .B2(new_n552), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n549), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT89), .Z(new_n684));
  NAND3_X1  g0484(.A1(new_n581), .A2(new_n590), .A3(new_n678), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  INV_X1    g0486(.A(new_n678), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n574), .B2(new_n580), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n596), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(G330), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT91), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n549), .A2(new_n678), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n591), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n687), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n215), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n463), .A2(G116), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n698), .A2(new_n253), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n223), .B2(new_n698), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n704));
  AND4_X1   g0504(.A1(new_n574), .A2(new_n580), .A3(new_n594), .A4(new_n592), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n636), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n591), .A2(new_n549), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n649), .A3(new_n643), .A4(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n657), .A2(new_n655), .A3(new_n649), .A4(new_n651), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n704), .A2(new_n708), .A3(new_n643), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n687), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n678), .B1(new_n659), .B2(new_n650), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n711), .B(new_n712), .C1(KEYINPUT29), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n637), .A2(new_n514), .A3(new_n553), .A4(new_n687), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n504), .A2(new_n593), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n544), .A2(new_n442), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n632), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n504), .A3(new_n593), .A4(new_n632), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n504), .A2(G179), .A3(new_n539), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n632), .B1(new_n527), .B2(new_n593), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n720), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n678), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n721), .A2(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n687), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n717), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  OAI21_X1  g0537(.A(new_n703), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(G13), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n247), .A3(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n253), .B1(new_n740), .B2(KEYINPUT94), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(KEYINPUT94), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n698), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n684), .B2(G330), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n684), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n251), .A3(KEYINPUT95), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G13), .B2(G33), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n683), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n743), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n215), .A2(G355), .A3(new_n261), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n697), .A2(new_n495), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n222), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n243), .A2(new_n247), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n754), .B1(G116), .B2(new_n215), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n218), .B1(G20), .B2(new_n340), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n753), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n219), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n266), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n219), .A2(G179), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G159), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n219), .A2(new_n442), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n765), .B(new_n771), .C1(G68), .C2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(G190), .A3(new_n378), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n767), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n355), .B1(new_n777), .B2(new_n292), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n773), .A2(new_n314), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n261), .B1(new_n781), .B2(new_n202), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G87), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n766), .A2(new_n314), .A3(G200), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n438), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n779), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n536), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT97), .Z(new_n791));
  INV_X1    g0591(.A(new_n777), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G311), .A2(new_n792), .B1(new_n769), .B2(G329), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n794), .B2(new_n776), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n780), .A2(G326), .ZN(new_n796));
  INV_X1    g0596(.A(new_n774), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n764), .A2(new_n800), .B1(new_n786), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n795), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n775), .A2(new_n788), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n752), .B(new_n761), .C1(new_n762), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n745), .A2(new_n805), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n444), .A2(new_n687), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n447), .A2(new_n450), .B1(new_n433), .B2(new_n678), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n444), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n714), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n809), .B(KEYINPUT99), .Z(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n714), .ZN(new_n813));
  INV_X1    g0613(.A(new_n735), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n743), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n780), .A2(G303), .B1(new_n792), .B2(G116), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n801), .B2(new_n797), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n536), .B1(new_n768), .B2(new_n821), .C1(new_n776), .C2(new_n800), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n765), .B1(G107), .B2(new_n784), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n462), .B2(new_n786), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n776), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G143), .B1(new_n792), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n781), .B2(new_n828), .C1(new_n829), .C2(new_n797), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n495), .B1(new_n834), .B2(new_n768), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n786), .A2(new_n239), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n202), .B2(new_n783), .C1(new_n355), .C2(new_n764), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n825), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n759), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n749), .A2(new_n759), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n753), .B1(new_n292), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n749), .B2(new_n809), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n817), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n602), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n220), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  OR3_X1    g0652(.A1(new_n222), .A2(new_n292), .A3(new_n356), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n253), .B(G13), .C1(new_n853), .C2(new_n238), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n364), .A2(new_n295), .ZN(new_n858));
  INV_X1    g0658(.A(new_n343), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT7), .B1(new_n495), .B2(G20), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n361), .A2(new_n348), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(G68), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n358), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n374), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT100), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n339), .B(new_n676), .C1(new_n340), .C2(new_n341), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT100), .B(new_n374), .C1(new_n858), .C2(new_n863), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n379), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n870), .A2(new_n365), .A3(new_n374), .A4(new_n386), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n857), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n867), .A2(new_n375), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n871), .A3(new_n857), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n676), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n866), .A2(new_n877), .A3(new_n868), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n664), .B2(new_n668), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n856), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  INV_X1    g0681(.A(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n389), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(KEYINPUT38), .C1(new_n872), .C2(new_n875), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT101), .B(new_n856), .C1(new_n876), .C2(new_n879), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n313), .A2(new_n678), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n676), .B1(new_n365), .B2(new_n374), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n389), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(new_n389), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n387), .A2(new_n375), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT102), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n857), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n873), .A2(new_n871), .A3(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(KEYINPUT103), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n874), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n895), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n884), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n888), .A2(new_n889), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n668), .A2(new_n877), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n885), .A2(new_n886), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n312), .A2(new_n678), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n313), .A2(new_n318), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n312), .B(new_n678), .C1(new_n287), .C2(new_n662), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n811), .B2(new_n807), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n909), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n454), .B1(new_n713), .B2(new_n715), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n671), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n732), .B2(KEYINPUT31), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n729), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n717), .A2(new_n923), .A3(new_n924), .A4(new_n733), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n809), .B1(new_n912), .B2(new_n913), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(new_n885), .A3(new_n929), .A4(new_n886), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n389), .A2(new_n892), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT104), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n389), .A2(new_n891), .A3(new_n892), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n898), .A2(KEYINPUT103), .A3(new_n899), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT103), .B1(new_n898), .B2(new_n899), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n935), .A2(new_n936), .A3(new_n875), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n856), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n927), .B1(new_n938), .B2(new_n884), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n930), .B1(new_n939), .B2(new_n929), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n455), .A2(new_n925), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  INV_X1    g0743(.A(G330), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n921), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(G1), .B1(new_n739), .B2(G20), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n921), .B2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n855), .B1(new_n946), .B2(new_n948), .ZN(G367));
  AOI21_X1  g0749(.A(new_n687), .B1(new_n604), .B2(new_n608), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n636), .A2(new_n950), .B1(new_n628), .B2(new_n687), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n693), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT42), .Z(new_n953));
  XOR2_X1   g0753(.A(new_n951), .B(KEYINPUT106), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n628), .B1(new_n954), .B2(new_n591), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n687), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n484), .A2(new_n687), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n644), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n643), .A2(new_n649), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n957), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n953), .A2(new_n956), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n961), .B(new_n962), .Z(new_n963));
  OR2_X1    g0763(.A1(new_n691), .A2(new_n954), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT107), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT107), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n963), .A2(new_n964), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n742), .B(KEYINPUT109), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n695), .A2(new_n951), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n695), .A2(new_n951), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n691), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n684), .A2(G330), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n689), .A2(new_n692), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n693), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n737), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n737), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n698), .B(KEYINPUT41), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n971), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n969), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n755), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n233), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n760), .B1(new_n215), .B2(new_n430), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n743), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G159), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n797), .A2(new_n993), .B1(new_n786), .B2(new_n292), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G58), .B2(new_n784), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n776), .A2(new_n829), .B1(new_n777), .B2(new_n202), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n536), .B(new_n996), .C1(G137), .C2(new_n769), .ZN(new_n997));
  INV_X1    g0797(.A(new_n764), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G68), .A2(new_n998), .B1(new_n780), .B2(G143), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n781), .A2(new_n821), .B1(new_n438), .B2(new_n764), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G294), .B2(new_n774), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n776), .A2(new_n789), .B1(new_n777), .B2(new_n801), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G317), .B2(new_n769), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n786), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n495), .B1(G97), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n783), .A2(new_n516), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n992), .B1(new_n1012), .B2(new_n759), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n751), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n960), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n988), .A2(new_n1016), .ZN(G387));
  INV_X1    g0817(.A(new_n698), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n983), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n737), .B2(new_n982), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n689), .A2(new_n1014), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n755), .B1(new_n229), .B2(new_n247), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n215), .A2(new_n261), .A3(new_n700), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n366), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT50), .B1(new_n366), .B2(G50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n699), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1024), .A2(new_n1028), .B1(new_n438), .B2(new_n697), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n760), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n743), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n776), .A2(new_n202), .B1(new_n777), .B2(new_n239), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G150), .B2(new_n769), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n429), .A2(new_n998), .B1(new_n780), .B2(G159), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n774), .A2(new_n408), .B1(new_n784), .B2(G77), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n611), .B1(G97), .B2(new_n1005), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n495), .B1(G326), .B2(new_n769), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n826), .A2(G317), .B1(new_n792), .B2(G303), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n781), .B2(new_n794), .C1(new_n821), .C2(new_n797), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n998), .A2(G283), .B1(new_n784), .B2(G294), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT49), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT111), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1038), .B1(new_n516), .B2(new_n786), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1046), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(KEYINPUT111), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1037), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1031), .B1(new_n1051), .B2(new_n759), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n982), .A2(new_n970), .B1(new_n1021), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1020), .A2(new_n1053), .ZN(G393));
  OR3_X1    g0854(.A1(new_n978), .A2(new_n983), .A3(KEYINPUT114), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT114), .B1(new_n978), .B2(new_n983), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n698), .A3(new_n984), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n780), .B1(new_n826), .B2(G311), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n536), .B1(new_n777), .B2(new_n800), .C1(new_n438), .C2(new_n786), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n797), .A2(new_n789), .B1(new_n516), .B2(new_n764), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n783), .A2(new_n801), .B1(new_n768), .B2(new_n794), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT113), .Z(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n780), .B1(new_n826), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n764), .A2(new_n292), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G50), .B2(new_n774), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n408), .A2(new_n792), .B1(new_n769), .B2(G143), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n784), .A2(G68), .B1(new_n1005), .B2(G87), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n495), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1063), .A2(new_n1065), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n759), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n989), .A2(new_n237), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n760), .B1(new_n266), .B2(new_n215), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n743), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1074), .B(new_n1077), .C1(new_n954), .C2(new_n751), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n978), .A2(KEYINPUT112), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n971), .B1(new_n978), .B2(KEYINPUT112), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1081), .ZN(G390));
  AOI21_X1  g0882(.A(KEYINPUT39), .B1(new_n938), .B2(new_n884), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n750), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n842), .A2(new_n366), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n797), .A2(new_n438), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1068), .B(new_n1088), .C1(G283), .C2(new_n780), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n776), .A2(new_n516), .B1(new_n768), .B2(new_n800), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n261), .B(new_n1090), .C1(G97), .C2(new_n792), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n785), .A3(new_n837), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n781), .A2(new_n1093), .B1(new_n786), .B2(new_n202), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n797), .A2(new_n828), .B1(new_n993), .B2(new_n764), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n783), .A2(new_n829), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1097), .B(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n536), .B1(new_n792), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n826), .A2(G132), .B1(new_n769), .B2(G125), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1096), .A2(new_n1099), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1092), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n743), .B(new_n1087), .C1(new_n1105), .C2(new_n762), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1086), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n889), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n807), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n714), .B2(new_n810), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n915), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n808), .A2(new_n444), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n710), .A2(new_n687), .A3(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1114), .A2(new_n807), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1108), .B1(new_n905), .B2(new_n906), .C1(new_n1115), .C2(new_n915), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n735), .A2(new_n810), .A3(new_n914), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n904), .A2(new_n933), .A3(new_n932), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n906), .B1(new_n1119), .B2(new_n856), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n915), .B1(new_n1114), .B2(new_n807), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n889), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n888), .A2(new_n907), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n1111), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n925), .A2(new_n926), .A3(G330), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT115), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT115), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n925), .A2(new_n926), .A3(new_n1127), .A4(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(KEYINPUT116), .B(new_n1118), .C1(new_n1124), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT116), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1129), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1107), .B1(new_n1135), .B2(new_n970), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n925), .A2(G330), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n454), .A2(new_n1137), .ZN(new_n1138));
  OR3_X1    g0938(.A1(new_n919), .A2(new_n671), .A3(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1117), .A2(new_n1115), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n812), .A2(G330), .A3(new_n925), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n915), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1110), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n734), .A2(new_n810), .A3(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n915), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1126), .A2(new_n1128), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1140), .A2(new_n1142), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1139), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n698), .B1(new_n1135), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(KEYINPUT116), .B(new_n1130), .C1(new_n1112), .C2(new_n1116), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1133), .B1(new_n1132), .B2(new_n1129), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1136), .B1(new_n1149), .B2(new_n1154), .ZN(G378));
  NOR3_X1   g0955(.A1(new_n919), .A2(new_n671), .A3(new_n1138), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n419), .A2(new_n425), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n422), .A3(new_n877), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n422), .A2(new_n877), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n419), .A2(new_n425), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT120), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1165), .A3(new_n1161), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1164), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n909), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n678), .B(new_n809), .C1(new_n659), .C2(new_n650), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n914), .B1(new_n1172), .B2(new_n1109), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1173), .B2(new_n887), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1085), .B2(new_n889), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n940), .A2(G330), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT40), .B1(new_n1120), .B2(new_n927), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n944), .B1(new_n1178), .B2(new_n930), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n918), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1170), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n918), .A2(new_n1179), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n1169), .A3(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1157), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1139), .B1(new_n1135), .B2(new_n1148), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n698), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1169), .A2(new_n750), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n495), .A2(G41), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G50), .B(new_n1192), .C1(new_n251), .C2(new_n246), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n781), .A2(new_n516), .B1(new_n786), .B2(new_n355), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G97), .B2(new_n774), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n776), .A2(new_n438), .B1(new_n768), .B2(new_n801), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n429), .B2(new_n792), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n998), .A2(G68), .B1(new_n784), .B2(G77), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1192), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n826), .A2(G128), .B1(new_n792), .B2(G137), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n783), .B2(new_n1100), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G150), .A2(new_n998), .B1(new_n780), .B2(G125), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT118), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G132), .C2(new_n774), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n993), .B2(new_n786), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1201), .B1(new_n1200), .B2(new_n1199), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n759), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n753), .B1(new_n202), .B2(new_n842), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1191), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1185), .B2(new_n970), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1190), .A2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n1146), .A2(new_n1143), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1142), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n970), .B(KEYINPUT121), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n915), .A2(new_n749), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n749), .A2(new_n759), .A3(G68), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n797), .A2(new_n516), .B1(new_n781), .B2(new_n800), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G97), .B2(new_n784), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n776), .A2(new_n801), .B1(new_n777), .B2(new_n438), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n261), .B(new_n1228), .C1(G303), .C2(new_n769), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n998), .A2(new_n429), .B1(new_n1005), .B2(G77), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT122), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n777), .A2(new_n829), .B1(new_n768), .B2(new_n1093), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G137), .B2(new_n826), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G50), .A2(new_n998), .B1(new_n780), .B2(G132), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n774), .A2(new_n1101), .B1(new_n784), .B2(G159), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n611), .B1(G58), .B2(new_n1005), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1233), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n753), .B(new_n1225), .C1(new_n1241), .C2(new_n759), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1222), .A2(new_n1223), .B1(new_n1224), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1148), .A2(new_n986), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1156), .A2(new_n1222), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(G381));
  NOR4_X1   g1046(.A1(G387), .A2(G390), .A3(G378), .A4(G381), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n846), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT123), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1190), .A3(new_n1218), .A4(new_n1250), .ZN(G407));
  INV_X1    g1051(.A(new_n1107), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1152), .B2(new_n971), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1135), .A2(new_n1148), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1018), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n677), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  INV_X1    g1059(.A(G213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(G343), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1218), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1187), .A2(new_n986), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1223), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1263), .A2(new_n1265), .B1(new_n1191), .B2(new_n1216), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1256), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1261), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1156), .B2(new_n1222), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1018), .B1(new_n1156), .B2(new_n1222), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1243), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n846), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(G384), .A3(new_n1243), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT124), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(G2897), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1273), .A2(G384), .A3(new_n1243), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1273), .B2(new_n1243), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1281), .B(new_n1280), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1279), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1259), .B1(new_n1268), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT125), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1290), .B(new_n1259), .C1(new_n1268), .C2(new_n1287), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1262), .A2(new_n1267), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1261), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1278), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1291), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1268), .A2(KEYINPUT62), .A3(new_n1278), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1278), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT127), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1297), .A2(new_n1291), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1299), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .A4(new_n1289), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1020), .A2(new_n1053), .B1(new_n805), .B2(new_n745), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1248), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(G390), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1058), .B(new_n1081), .C1(new_n1248), .C2(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(G387), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1303), .A2(new_n1308), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G387), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1313), .B(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1288), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1294), .B(KEYINPUT63), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1277), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1277), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1314), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1323), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1317), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(G402));
endmodule


