

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774;

  AND2_X1 U371 ( .A1(n764), .A2(n640), .ZN(n391) );
  INV_X2 U372 ( .A(G146), .ZN(n462) );
  XNOR2_X2 U373 ( .A(n428), .B(n604), .ZN(n714) );
  XOR2_X2 U374 ( .A(KEYINPUT89), .B(KEYINPUT0), .Z(n396) );
  AND2_X2 U375 ( .A1(n653), .A2(KEYINPUT44), .ZN(n559) );
  XNOR2_X1 U376 ( .A(G143), .B(G113), .ZN(n501) );
  XOR2_X1 U377 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n757) );
  AND2_X2 U378 ( .A1(n454), .A2(KEYINPUT67), .ZN(n424) );
  NAND2_X2 U379 ( .A1(n470), .A2(n469), .ZN(n382) );
  AND2_X1 U380 ( .A1(n456), .A2(n467), .ZN(n455) );
  INV_X2 U381 ( .A(n676), .ZN(n349) );
  XNOR2_X1 U382 ( .A(G107), .B(G104), .ZN(n411) );
  NAND2_X1 U383 ( .A1(n453), .A2(n455), .ZN(n470) );
  NAND2_X1 U384 ( .A1(n745), .A2(n451), .ZN(n646) );
  AND2_X1 U385 ( .A1(n764), .A2(n645), .ZN(n451) );
  XNOR2_X1 U386 ( .A(n408), .B(KEYINPUT35), .ZN(n581) );
  AND2_X1 U387 ( .A1(n717), .A2(n606), .ZN(n596) );
  XNOR2_X1 U388 ( .A(n487), .B(KEYINPUT19), .ZN(n611) );
  XNOR2_X1 U389 ( .A(n411), .B(n410), .ZN(n740) );
  INV_X1 U390 ( .A(KEYINPUT8), .ZN(n378) );
  INV_X1 U391 ( .A(KEYINPUT60), .ZN(n357) );
  INV_X1 U392 ( .A(KEYINPUT56), .ZN(n350) );
  NAND2_X1 U393 ( .A1(n424), .A2(n468), .ZN(n453) );
  NAND2_X1 U394 ( .A1(n365), .A2(n418), .ZN(n364) );
  NAND2_X1 U395 ( .A1(n395), .A2(n368), .ZN(n367) );
  NAND2_X1 U396 ( .A1(n583), .A2(KEYINPUT86), .ZN(n368) );
  NAND2_X1 U397 ( .A1(n617), .A2(n441), .ZN(n465) );
  AND2_X1 U398 ( .A1(n389), .A2(n442), .ZN(n441) );
  NAND2_X1 U399 ( .A1(n555), .A2(n608), .ZN(n408) );
  INV_X1 U400 ( .A(n682), .ZN(n433) );
  NAND2_X1 U401 ( .A1(n466), .A2(n516), .ZN(n518) );
  NAND2_X1 U402 ( .A1(n552), .A2(n618), .ZN(n407) );
  XNOR2_X1 U403 ( .A(n375), .B(KEYINPUT95), .ZN(n606) );
  NAND2_X1 U404 ( .A1(n377), .A2(n376), .ZN(n375) );
  XNOR2_X1 U405 ( .A(n563), .B(KEYINPUT6), .ZN(n618) );
  INV_X1 U406 ( .A(n674), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n673), .B(n672), .ZN(n674) );
  OR2_X1 U408 ( .A1(n619), .A2(n597), .ZN(n700) );
  INV_X1 U409 ( .A(n661), .ZN(n361) );
  XNOR2_X1 U410 ( .A(n463), .B(n459), .ZN(n656) );
  XOR2_X1 U411 ( .A(KEYINPUT59), .B(n660), .Z(n661) );
  XNOR2_X1 U412 ( .A(n544), .B(n464), .ZN(n463) );
  XNOR2_X1 U413 ( .A(n753), .B(n460), .ZN(n459) );
  XNOR2_X1 U414 ( .A(n379), .B(n378), .ZN(n543) );
  XNOR2_X1 U415 ( .A(n520), .B(G137), .ZN(n452) );
  XNOR2_X1 U416 ( .A(n539), .B(n541), .ZN(n460) );
  NAND2_X1 U417 ( .A1(G237), .A2(G234), .ZN(n488) );
  XNOR2_X1 U418 ( .A(KEYINPUT77), .B(KEYINPUT17), .ZN(n479) );
  XNOR2_X1 U419 ( .A(KEYINPUT18), .B(KEYINPUT91), .ZN(n478) );
  XNOR2_X1 U420 ( .A(G122), .B(G104), .ZN(n500) );
  XOR2_X1 U421 ( .A(G140), .B(KEYINPUT93), .Z(n522) );
  XNOR2_X1 U422 ( .A(G140), .B(KEYINPUT10), .ZN(n461) );
  XNOR2_X2 U423 ( .A(n426), .B(n425), .ZN(n374) );
  XNOR2_X1 U424 ( .A(n351), .B(n350), .ZN(G51) );
  NAND2_X1 U425 ( .A1(n355), .A2(n349), .ZN(n351) );
  XNOR2_X1 U426 ( .A(n352), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U427 ( .A1(n353), .A2(n349), .ZN(n352) );
  XNOR2_X1 U428 ( .A(n650), .B(n354), .ZN(n353) );
  INV_X1 U429 ( .A(n649), .ZN(n354) );
  XNOR2_X1 U430 ( .A(n675), .B(n356), .ZN(n355) );
  XNOR2_X1 U431 ( .A(n358), .B(n357), .ZN(G60) );
  NAND2_X1 U432 ( .A1(n360), .A2(n349), .ZN(n358) );
  XNOR2_X1 U433 ( .A(n359), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U434 ( .A1(n362), .A2(n349), .ZN(n359) );
  XNOR2_X1 U435 ( .A(n662), .B(n361), .ZN(n360) );
  XNOR2_X2 U436 ( .A(n450), .B(n558), .ZN(n653) );
  XNOR2_X1 U437 ( .A(n413), .B(n481), .ZN(n412) );
  XNOR2_X1 U438 ( .A(n652), .B(n363), .ZN(n362) );
  INV_X1 U439 ( .A(n651), .ZN(n363) );
  NAND2_X1 U440 ( .A1(n370), .A2(KEYINPUT45), .ZN(n369) );
  NAND2_X1 U441 ( .A1(n423), .A2(n422), .ZN(n370) );
  NAND2_X2 U442 ( .A1(n366), .A2(n364), .ZN(n745) );
  INV_X1 U443 ( .A(n370), .ZN(n365) );
  AND2_X2 U444 ( .A1(n369), .A2(n367), .ZN(n366) );
  XNOR2_X2 U445 ( .A(n755), .B(n373), .ZN(n372) );
  XNOR2_X2 U446 ( .A(n371), .B(n526), .ZN(n601) );
  NAND2_X1 U447 ( .A1(n664), .A2(n545), .ZN(n371) );
  XNOR2_X2 U448 ( .A(n372), .B(n525), .ZN(n664) );
  INV_X1 U449 ( .A(n524), .ZN(n373) );
  NAND2_X1 U450 ( .A1(n374), .A2(G472), .ZN(n650) );
  NAND2_X1 U451 ( .A1(n374), .A2(G210), .ZN(n675) );
  INV_X1 U452 ( .A(n606), .ZN(n595) );
  INV_X1 U453 ( .A(n601), .ZN(n376) );
  INV_X1 U454 ( .A(n700), .ZN(n377) );
  NAND2_X1 U455 ( .A1(n543), .A2(G221), .ZN(n544) );
  NAND2_X1 U456 ( .A1(n766), .A2(G234), .ZN(n379) );
  INV_X4 U457 ( .A(G953), .ZN(n766) );
  BUF_X1 U458 ( .A(n437), .Z(n380) );
  BUF_X1 U459 ( .A(n528), .Z(n381) );
  BUF_X1 U460 ( .A(n692), .Z(n383) );
  NAND2_X1 U461 ( .A1(n470), .A2(n469), .ZN(n426) );
  NOR2_X1 U462 ( .A1(n611), .A2(n493), .ZN(n384) );
  NOR2_X1 U463 ( .A1(n611), .A2(n493), .ZN(n494) );
  BUF_X1 U464 ( .A(n745), .Z(n385) );
  XNOR2_X1 U465 ( .A(n384), .B(n396), .ZN(n386) );
  XNOR2_X1 U466 ( .A(n494), .B(n396), .ZN(n466) );
  XNOR2_X1 U467 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n517) );
  NAND2_X1 U468 ( .A1(n434), .A2(n433), .ZN(n630) );
  INV_X1 U469 ( .A(n721), .ZN(n434) );
  NOR2_X1 U470 ( .A1(n630), .A2(n431), .ZN(n443) );
  NAND2_X1 U471 ( .A1(n432), .A2(KEYINPUT80), .ZN(n431) );
  INV_X1 U472 ( .A(KEYINPUT47), .ZN(n432) );
  NAND2_X1 U473 ( .A1(n695), .A2(n629), .ZN(n444) );
  XNOR2_X1 U474 ( .A(n757), .B(n447), .ZN(n527) );
  XNOR2_X1 U475 ( .A(G101), .B(KEYINPUT70), .ZN(n447) );
  INV_X1 U476 ( .A(G237), .ZN(n483) );
  XOR2_X1 U477 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n531) );
  XNOR2_X1 U478 ( .A(n527), .B(G146), .ZN(n446) );
  NAND2_X1 U479 ( .A1(n583), .A2(n399), .ZN(n420) );
  NAND2_X1 U480 ( .A1(n770), .A2(n421), .ZN(n419) );
  XNOR2_X1 U481 ( .A(G119), .B(G116), .ZN(n473) );
  NOR2_X1 U482 ( .A1(G953), .A2(G237), .ZN(n529) );
  XNOR2_X1 U483 ( .A(n504), .B(G475), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n465), .B(n397), .ZN(n639) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n508) );
  XNOR2_X1 U486 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n506), .B(KEYINPUT103), .ZN(n430) );
  XNOR2_X1 U488 ( .A(G107), .B(KEYINPUT9), .ZN(n506) );
  XNOR2_X1 U489 ( .A(n405), .B(n390), .ZN(n404) );
  XNOR2_X1 U490 ( .A(n500), .B(n501), .ZN(n405) );
  XNOR2_X1 U491 ( .A(KEYINPUT11), .B(KEYINPUT97), .ZN(n498) );
  XOR2_X1 U492 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n499) );
  AND2_X1 U493 ( .A1(n701), .A2(n563), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n570) );
  XNOR2_X1 U495 ( .A(n512), .B(G478), .ZN(n435) );
  OR2_X1 U496 ( .A1(n651), .A2(G902), .ZN(n436) );
  INV_X1 U497 ( .A(KEYINPUT45), .ZN(n421) );
  XNOR2_X1 U498 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  XNOR2_X1 U499 ( .A(n409), .B(n605), .ZN(n617) );
  NOR2_X1 U500 ( .A1(n444), .A2(n443), .ZN(n442) );
  INV_X1 U501 ( .A(KEYINPUT66), .ZN(n425) );
  XNOR2_X1 U502 ( .A(n601), .B(KEYINPUT1), .ZN(n551) );
  INV_X1 U503 ( .A(G902), .ZN(n545) );
  XNOR2_X1 U504 ( .A(n535), .B(n534), .ZN(n648) );
  INV_X1 U505 ( .A(G110), .ZN(n410) );
  XNOR2_X1 U506 ( .A(KEYINPUT16), .B(G122), .ZN(n476) );
  XNOR2_X1 U507 ( .A(n540), .B(n542), .ZN(n464) );
  XNOR2_X1 U508 ( .A(n523), .B(G146), .ZN(n524) );
  NAND2_X1 U509 ( .A1(n618), .A2(n445), .ZN(n621) );
  AND2_X1 U510 ( .A1(n620), .A2(n393), .ZN(n445) );
  NOR2_X2 U511 ( .A1(n720), .A2(n719), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n458), .B(KEYINPUT39), .ZN(n636) );
  NAND2_X1 U513 ( .A1(n596), .A2(n607), .ZN(n458) );
  BUF_X1 U514 ( .A(n551), .Z(n701) );
  NAND2_X1 U515 ( .A1(n401), .A2(n570), .ZN(n622) );
  XOR2_X1 U516 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  XNOR2_X1 U517 ( .A(n511), .B(n510), .ZN(n651) );
  XNOR2_X1 U518 ( .A(G116), .B(G122), .ZN(n507) );
  XNOR2_X1 U519 ( .A(n503), .B(n403), .ZN(n660) );
  XNOR2_X1 U520 ( .A(n753), .B(n497), .ZN(n503) );
  XNOR2_X1 U521 ( .A(n502), .B(n404), .ZN(n403) );
  NOR2_X1 U522 ( .A1(n766), .A2(G952), .ZN(n676) );
  INV_X1 U523 ( .A(KEYINPUT109), .ZN(n472) );
  INV_X1 U524 ( .A(n622), .ZN(n689) );
  XNOR2_X1 U525 ( .A(n505), .B(n402), .ZN(n569) );
  INV_X1 U526 ( .A(n569), .ZN(n401) );
  BUF_X1 U527 ( .A(n581), .Z(n770) );
  AND2_X1 U528 ( .A1(n546), .A2(G217), .ZN(n387) );
  OR2_X1 U529 ( .A1(n595), .A2(n707), .ZN(n388) );
  AND2_X1 U530 ( .A1(n616), .A2(n615), .ZN(n389) );
  XNOR2_X1 U531 ( .A(KEYINPUT100), .B(KEYINPUT98), .ZN(n390) );
  AND2_X1 U532 ( .A1(n560), .A2(n559), .ZN(n392) );
  AND2_X1 U533 ( .A1(n716), .A2(n619), .ZN(n393) );
  NOR2_X1 U534 ( .A1(n557), .A2(n701), .ZN(n394) );
  AND2_X1 U535 ( .A1(n584), .A2(KEYINPUT45), .ZN(n395) );
  XNOR2_X1 U536 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n397) );
  AND2_X1 U537 ( .A1(n645), .A2(n471), .ZN(n398) );
  AND2_X1 U538 ( .A1(n421), .A2(KEYINPUT86), .ZN(n399) );
  AND2_X1 U539 ( .A1(n471), .A2(KEYINPUT83), .ZN(n400) );
  INV_X1 U540 ( .A(KEYINPUT67), .ZN(n471) );
  NAND2_X1 U541 ( .A1(n406), .A2(G478), .ZN(n652) );
  XNOR2_X1 U542 ( .A(n755), .B(n446), .ZN(n535) );
  XNOR2_X2 U543 ( .A(n382), .B(n425), .ZN(n406) );
  XNOR2_X2 U544 ( .A(n407), .B(KEYINPUT33), .ZN(n698) );
  NAND2_X1 U545 ( .A1(n647), .A2(KEYINPUT2), .ZN(n469) );
  NAND2_X1 U546 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U547 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U548 ( .A1(n772), .A2(n773), .ZN(n409) );
  XNOR2_X2 U549 ( .A(n635), .B(n594), .ZN(n717) );
  AND2_X1 U550 ( .A1(n580), .A2(n579), .ZN(n422) );
  AND2_X1 U551 ( .A1(n556), .A2(n701), .ZN(n576) );
  XNOR2_X1 U552 ( .A(n741), .B(n412), .ZN(n449) );
  XNOR2_X1 U553 ( .A(n415), .B(n414), .ZN(n413) );
  XNOR2_X2 U554 ( .A(n528), .B(n476), .ZN(n741) );
  XNOR2_X2 U555 ( .A(n416), .B(n473), .ZN(n528) );
  XNOR2_X1 U556 ( .A(n479), .B(n477), .ZN(n414) );
  XNOR2_X1 U557 ( .A(n417), .B(n480), .ZN(n415) );
  XNOR2_X2 U558 ( .A(n475), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U559 ( .A(n417), .B(G134), .ZN(n519) );
  XNOR2_X2 U560 ( .A(G143), .B(G128), .ZN(n417) );
  NAND2_X1 U561 ( .A1(n562), .A2(n561), .ZN(n423) );
  XNOR2_X1 U562 ( .A(n440), .B(n538), .ZN(n439) );
  XNOR2_X2 U563 ( .A(n427), .B(KEYINPUT42), .ZN(n772) );
  NAND2_X1 U564 ( .A1(n714), .A2(n614), .ZN(n427) );
  NAND2_X1 U565 ( .A1(n392), .A2(n437), .ZN(n562) );
  NAND2_X1 U566 ( .A1(n437), .A2(n474), .ZN(n583) );
  XNOR2_X1 U567 ( .A(n380), .B(G110), .ZN(G12) );
  XNOR2_X2 U568 ( .A(n550), .B(n472), .ZN(n437) );
  NAND2_X1 U569 ( .A1(n556), .A2(n438), .ZN(n440) );
  NAND2_X1 U570 ( .A1(n439), .A2(n619), .ZN(n550) );
  AND2_X1 U571 ( .A1(n385), .A2(n764), .ZN(n647) );
  XNOR2_X2 U572 ( .A(n448), .B(n484), .ZN(n593) );
  NAND2_X1 U573 ( .A1(n670), .A2(n643), .ZN(n448) );
  XNOR2_X1 U574 ( .A(n449), .B(n525), .ZN(n670) );
  NAND2_X1 U575 ( .A1(n556), .A2(n394), .ZN(n450) );
  NAND2_X1 U576 ( .A1(n745), .A2(n391), .ZN(n642) );
  XNOR2_X2 U577 ( .A(n519), .B(n452), .ZN(n755) );
  NAND2_X1 U578 ( .A1(n646), .A2(KEYINPUT83), .ZN(n454) );
  NAND2_X1 U579 ( .A1(n644), .A2(n398), .ZN(n456) );
  XNOR2_X2 U580 ( .A(n457), .B(KEYINPUT40), .ZN(n773) );
  NAND2_X1 U581 ( .A1(n636), .A2(n689), .ZN(n457) );
  XNOR2_X2 U582 ( .A(n495), .B(n461), .ZN(n753) );
  XNOR2_X2 U583 ( .A(n462), .B(G125), .ZN(n495) );
  INV_X1 U584 ( .A(n386), .ZN(n566) );
  NOR2_X1 U585 ( .A1(n566), .A2(n388), .ZN(n678) );
  NAND2_X1 U586 ( .A1(n698), .A2(n386), .ZN(n554) );
  NAND2_X1 U587 ( .A1(n646), .A2(n400), .ZN(n467) );
  NAND2_X1 U588 ( .A1(n644), .A2(n645), .ZN(n468) );
  AND2_X1 U589 ( .A1(n653), .A2(n582), .ZN(n474) );
  INV_X1 U590 ( .A(KEYINPUT24), .ZN(n541) );
  BUF_X1 U591 ( .A(n698), .Z(n724) );
  XNOR2_X1 U592 ( .A(n533), .B(n532), .ZN(n534) );
  BUF_X1 U593 ( .A(n670), .Z(n673) );
  XNOR2_X2 U594 ( .A(G113), .B(KEYINPUT72), .ZN(n475) );
  NAND2_X1 U595 ( .A1(G224), .A2(n766), .ZN(n477) );
  INV_X1 U596 ( .A(n478), .ZN(n480) );
  XOR2_X1 U597 ( .A(n495), .B(KEYINPUT90), .Z(n481) );
  XNOR2_X1 U598 ( .A(n740), .B(KEYINPUT73), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n527), .B(n482), .ZN(n525) );
  NAND2_X1 U600 ( .A1(n545), .A2(n483), .ZN(n485) );
  NAND2_X1 U601 ( .A1(n485), .A2(G210), .ZN(n484) );
  NAND2_X1 U602 ( .A1(n485), .A2(G214), .ZN(n716) );
  INV_X1 U603 ( .A(n716), .ZN(n486) );
  NOR2_X2 U604 ( .A1(n593), .A2(n486), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n488), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U606 ( .A1(n491), .A2(G902), .ZN(n489) );
  XOR2_X1 U607 ( .A(KEYINPUT92), .B(n489), .Z(n490) );
  NAND2_X1 U608 ( .A1(G953), .A2(n490), .ZN(n587) );
  NOR2_X1 U609 ( .A1(n587), .A2(G898), .ZN(n492) );
  NAND2_X1 U610 ( .A1(G952), .A2(n491), .ZN(n732) );
  NOR2_X1 U611 ( .A1(n732), .A2(G953), .ZN(n590) );
  NOR2_X1 U612 ( .A1(n492), .A2(n590), .ZN(n493) );
  NAND2_X1 U613 ( .A1(n529), .A2(G214), .ZN(n496) );
  XNOR2_X2 U614 ( .A(KEYINPUT71), .B(G131), .ZN(n520) );
  XNOR2_X1 U615 ( .A(n496), .B(n520), .ZN(n497) );
  XNOR2_X1 U616 ( .A(n499), .B(n498), .ZN(n502) );
  NOR2_X1 U617 ( .A1(G902), .A2(n660), .ZN(n505) );
  XNOR2_X1 U618 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n504) );
  XNOR2_X1 U619 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U620 ( .A(n508), .B(n507), .ZN(n511) );
  AND2_X1 U621 ( .A1(n543), .A2(G217), .ZN(n509) );
  XNOR2_X1 U622 ( .A(n519), .B(n509), .ZN(n510) );
  NAND2_X1 U623 ( .A1(n569), .A2(n570), .ZN(n719) );
  NAND2_X1 U624 ( .A1(n643), .A2(G234), .ZN(n513) );
  XNOR2_X1 U625 ( .A(n513), .B(KEYINPUT20), .ZN(n546) );
  AND2_X1 U626 ( .A1(n546), .A2(G221), .ZN(n515) );
  INV_X1 U627 ( .A(KEYINPUT21), .ZN(n514) );
  XNOR2_X1 U628 ( .A(n515), .B(n514), .ZN(n597) );
  NOR2_X1 U629 ( .A1(n719), .A2(n597), .ZN(n516) );
  XNOR2_X2 U630 ( .A(n518), .B(n517), .ZN(n556) );
  NAND2_X1 U631 ( .A1(G227), .A2(n766), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U633 ( .A(G469), .ZN(n526) );
  INV_X1 U634 ( .A(n381), .ZN(n533) );
  NAND2_X1 U635 ( .A1(n529), .A2(G210), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U637 ( .A1(n648), .A2(n545), .ZN(n537) );
  INV_X1 U638 ( .A(G472), .ZN(n536) );
  XNOR2_X2 U639 ( .A(n537), .B(n536), .ZN(n563) );
  INV_X1 U640 ( .A(KEYINPUT68), .ZN(n538) );
  XOR2_X1 U641 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n540) );
  XNOR2_X1 U642 ( .A(G137), .B(G110), .ZN(n539) );
  XNOR2_X1 U643 ( .A(G128), .B(G119), .ZN(n542) );
  NAND2_X1 U644 ( .A1(n656), .A2(n545), .ZN(n549) );
  XOR2_X1 U645 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n547) );
  XNOR2_X1 U646 ( .A(n547), .B(n387), .ZN(n548) );
  XNOR2_X2 U647 ( .A(n549), .B(n548), .ZN(n619) );
  NOR2_X2 U648 ( .A1(n551), .A2(n700), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n564), .B(KEYINPUT110), .ZN(n552) );
  XOR2_X1 U650 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n553) );
  XNOR2_X1 U651 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U652 ( .A1(n570), .A2(n569), .ZN(n608) );
  NAND2_X1 U653 ( .A1(n581), .A2(KEYINPUT86), .ZN(n560) );
  XNOR2_X1 U654 ( .A(n619), .B(KEYINPUT107), .ZN(n703) );
  OR2_X1 U655 ( .A1(n618), .A2(n703), .ZN(n557) );
  XNOR2_X1 U656 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n558) );
  INV_X1 U657 ( .A(KEYINPUT44), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n582), .A2(KEYINPUT86), .ZN(n561) );
  INV_X1 U659 ( .A(n563), .ZN(n585) );
  BUF_X1 U660 ( .A(n585), .Z(n707) );
  NAND2_X1 U661 ( .A1(n564), .A2(n707), .ZN(n565) );
  XNOR2_X1 U662 ( .A(n565), .B(KEYINPUT96), .ZN(n711) );
  NOR2_X1 U663 ( .A1(n711), .A2(n566), .ZN(n568) );
  INV_X1 U664 ( .A(KEYINPUT31), .ZN(n567) );
  XNOR2_X1 U665 ( .A(n568), .B(n567), .ZN(n692) );
  OR2_X1 U666 ( .A1(n692), .A2(n678), .ZN(n572) );
  NOR2_X1 U667 ( .A1(n401), .A2(n570), .ZN(n691) );
  NOR2_X1 U668 ( .A1(n689), .A2(n691), .ZN(n721) );
  XOR2_X1 U669 ( .A(n721), .B(KEYINPUT80), .Z(n571) );
  NAND2_X1 U670 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U671 ( .A(n573), .B(KEYINPUT106), .ZN(n580) );
  INV_X1 U672 ( .A(n703), .ZN(n574) );
  NOR2_X1 U673 ( .A1(n618), .A2(n574), .ZN(n575) );
  NAND2_X1 U674 ( .A1(n576), .A2(n575), .ZN(n578) );
  INV_X1 U675 ( .A(KEYINPUT108), .ZN(n577) );
  XNOR2_X1 U676 ( .A(n578), .B(n577), .ZN(n774) );
  INV_X1 U677 ( .A(n774), .ZN(n579) );
  INV_X1 U678 ( .A(n770), .ZN(n584) );
  NAND2_X1 U679 ( .A1(n585), .A2(n716), .ZN(n586) );
  XOR2_X1 U680 ( .A(n586), .B(KEYINPUT30), .Z(n592) );
  NOR2_X1 U681 ( .A1(G900), .A2(n587), .ZN(n588) );
  XOR2_X1 U682 ( .A(KEYINPUT111), .B(n588), .Z(n589) );
  NOR2_X1 U683 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U684 ( .A(KEYINPUT79), .B(n591), .ZN(n598) );
  AND2_X1 U685 ( .A1(n592), .A2(n598), .ZN(n607) );
  BUF_X2 U686 ( .A(n593), .Z(n635) );
  XOR2_X1 U687 ( .A(KEYINPUT75), .B(KEYINPUT38), .Z(n594) );
  INV_X1 U688 ( .A(n597), .ZN(n704) );
  AND2_X1 U689 ( .A1(n598), .A2(n704), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n599) );
  NOR2_X1 U691 ( .A1(n563), .A2(n599), .ZN(n600) );
  XOR2_X1 U692 ( .A(KEYINPUT28), .B(n600), .Z(n603) );
  BUF_X1 U693 ( .A(n601), .Z(n602) );
  NOR2_X1 U694 ( .A1(n603), .A2(n602), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n717), .A2(n716), .ZN(n720) );
  XNOR2_X1 U696 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n604) );
  XOR2_X1 U697 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n605) );
  AND2_X1 U698 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U699 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U700 ( .A1(n610), .A2(n635), .ZN(n655) );
  XNOR2_X1 U701 ( .A(n655), .B(KEYINPUT81), .ZN(n616) );
  BUF_X1 U702 ( .A(n611), .Z(n612) );
  INV_X1 U703 ( .A(n612), .ZN(n613) );
  NAND2_X1 U704 ( .A1(n614), .A2(n613), .ZN(n682) );
  NAND2_X1 U705 ( .A1(KEYINPUT47), .A2(n630), .ZN(n615) );
  NOR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n631) );
  INV_X1 U707 ( .A(n635), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n631), .A2(n623), .ZN(n625) );
  XNOR2_X1 U709 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n624) );
  XNOR2_X1 U710 ( .A(n625), .B(n624), .ZN(n627) );
  INV_X1 U711 ( .A(n701), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n695) );
  NOR2_X1 U713 ( .A1(n682), .A2(KEYINPUT80), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n721), .A2(n628), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n631), .A2(n701), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(KEYINPUT112), .ZN(n633) );
  XNOR2_X1 U717 ( .A(n633), .B(KEYINPUT43), .ZN(n634) );
  AND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n636), .A2(n691), .ZN(n696) );
  INV_X1 U720 ( .A(n696), .ZN(n637) );
  NOR2_X1 U721 ( .A1(n654), .A2(n637), .ZN(n638) );
  AND2_X2 U722 ( .A1(n639), .A2(n638), .ZN(n764) );
  INV_X1 U723 ( .A(KEYINPUT83), .ZN(n640) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n641) );
  INV_X1 U725 ( .A(n643), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n653), .B(G119), .ZN(G21) );
  XOR2_X1 U727 ( .A(n654), .B(G140), .Z(G42) );
  XOR2_X1 U728 ( .A(G143), .B(n655), .Z(G45) );
  BUF_X1 U729 ( .A(n406), .Z(n663) );
  NAND2_X1 U730 ( .A1(n663), .A2(G217), .ZN(n658) );
  XOR2_X1 U731 ( .A(KEYINPUT122), .B(n656), .Z(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n659), .A2(n676), .ZN(G66) );
  NAND2_X1 U734 ( .A1(n406), .A2(G475), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n663), .A2(G469), .ZN(n668) );
  BUF_X1 U736 ( .A(n664), .Z(n666) );
  XNOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n669), .A2(n676), .ZN(G54) );
  XNOR2_X1 U741 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n671), .B(KEYINPUT55), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n678), .A2(n689), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(G104), .ZN(G6) );
  XOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n680) );
  NAND2_X1 U746 ( .A1(n678), .A2(n691), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(G107), .B(n681), .ZN(G9) );
  XOR2_X1 U749 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n684) );
  NAND2_X1 U750 ( .A1(n433), .A2(n691), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n686) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT114), .Z(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(G30) );
  NAND2_X1 U754 ( .A1(n433), .A2(n689), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(KEYINPUT116), .ZN(n688) );
  XNOR2_X1 U756 ( .A(G146), .B(n688), .ZN(G48) );
  NAND2_X1 U757 ( .A1(n383), .A2(n689), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(G113), .ZN(G15) );
  NAND2_X1 U759 ( .A1(n383), .A2(n691), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n693), .B(G116), .ZN(G18) );
  XOR2_X1 U761 ( .A(G125), .B(KEYINPUT37), .Z(n694) );
  XNOR2_X1 U762 ( .A(n695), .B(n694), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G134), .B(n696), .ZN(G36) );
  XNOR2_X1 U764 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n647), .B(n697), .ZN(n737) );
  NAND2_X1 U766 ( .A1(n714), .A2(n724), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n699), .B(KEYINPUT119), .ZN(n734) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U769 ( .A(KEYINPUT50), .B(n702), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U771 ( .A(KEYINPUT49), .B(n705), .Z(n706) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U775 ( .A(KEYINPUT51), .B(n712), .Z(n713) );
  NAND2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U777 ( .A(KEYINPUT117), .B(n715), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U781 ( .A1(n723), .A2(n722), .ZN(n726) );
  INV_X1 U782 ( .A(n724), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n727), .B(KEYINPUT118), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U786 ( .A(KEYINPUT52), .B(n730), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U789 ( .A(KEYINPUT120), .B(n735), .ZN(n736) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n738), .A2(G953), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n739), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U793 ( .A(n740), .B(G101), .Z(n742) );
  XNOR2_X1 U794 ( .A(n741), .B(n742), .ZN(n744) );
  NOR2_X1 U795 ( .A1(G898), .A2(n766), .ZN(n743) );
  NOR2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n752) );
  NAND2_X1 U797 ( .A1(n385), .A2(n766), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n747) );
  NAND2_X1 U799 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n747), .B(n746), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(G69) );
  XOR2_X1 U804 ( .A(KEYINPUT93), .B(n753), .Z(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n765) );
  INV_X1 U807 ( .A(n765), .ZN(n758) );
  XNOR2_X1 U808 ( .A(G227), .B(n758), .ZN(n759) );
  XNOR2_X1 U809 ( .A(n759), .B(KEYINPUT124), .ZN(n760) );
  NAND2_X1 U810 ( .A1(n760), .A2(G900), .ZN(n761) );
  XOR2_X1 U811 ( .A(KEYINPUT125), .B(n761), .Z(n762) );
  NAND2_X1 U812 ( .A1(G953), .A2(n762), .ZN(n763) );
  XNOR2_X1 U813 ( .A(KEYINPUT126), .B(n763), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n765), .B(n764), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G72) );
  XNOR2_X1 U817 ( .A(n770), .B(G122), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n771), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U819 ( .A(n772), .B(G137), .ZN(G39) );
  XNOR2_X1 U820 ( .A(n773), .B(G131), .ZN(G33) );
  XOR2_X1 U821 ( .A(G101), .B(n774), .Z(G3) );
endmodule

