//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  OR2_X1    g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  NOR2_X1   g0001(.A1(new_n201), .A2(G50), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AND2_X1   g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n201), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n210), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n213), .B1(new_n215), .B2(new_n216), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G274), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n246), .B1(new_n214), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n250), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(G226), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G223), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G222), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n262), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n254), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(G77), .C2(new_n262), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n257), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G200), .B2(new_n273), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G20), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n203), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n259), .A3(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G20), .B2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(G33), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n279), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n238), .B1(new_n249), .B2(G20), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(new_n295), .B1(new_n238), .B2(new_n293), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n291), .A2(KEYINPUT9), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n276), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n297), .B(new_n304), .C1(G179), .C2(new_n273), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n249), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n294), .A2(G77), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n309), .A2(new_n289), .B1(new_n280), .B2(new_n204), .ZN(new_n310));
  INV_X1    g0110(.A(new_n288), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n285), .ZN(new_n312));
  INV_X1    g0112(.A(new_n279), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n308), .B1(G77), .B2(new_n292), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n227), .B1(new_n260), .B2(new_n261), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT66), .B(G1698), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n315), .A2(new_n316), .B1(new_n319), .B2(G107), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n264), .B1(new_n260), .B2(new_n261), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n271), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n253), .B1(G244), .B2(new_n256), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n314), .B1(new_n328), .B2(G169), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(G179), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n274), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT68), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n314), .B1(G200), .B2(new_n327), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n306), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n319), .B2(new_n280), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n280), .A4(new_n261), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n282), .B2(new_n284), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n280), .B1(new_n201), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT72), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n285), .A2(G159), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n201), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n345), .A4(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n260), .A2(new_n280), .A3(new_n261), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n240), .B1(new_n355), .B2(new_n338), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n346), .A2(new_n349), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n351), .A2(new_n279), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n351), .A2(new_n358), .A3(KEYINPUT74), .A4(new_n279), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n294), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n311), .A2(new_n307), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n364), .A2(new_n365), .B1(new_n292), .B2(new_n311), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT18), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT75), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n265), .A2(new_n267), .A3(G223), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G226), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n319), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n372), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n316), .B2(G223), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT75), .B(new_n374), .C1(new_n378), .C2(new_n319), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n379), .A3(new_n271), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n252), .B1(new_n227), .B2(new_n255), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G169), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(G179), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n368), .A2(new_n369), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g0187(.A(KEYINPUT76), .B(G190), .Z(new_n388));
  NAND3_X1  g0188(.A1(new_n380), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n374), .B1(new_n378), .B2(new_n319), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n254), .B1(new_n390), .B2(new_n370), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n381), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(G200), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n363), .A2(new_n367), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n366), .B1(new_n361), .B2(new_n362), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n384), .A2(new_n385), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT18), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n393), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n387), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n286), .A2(new_n238), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n289), .A2(new_n204), .B1(new_n280), .B2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n279), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT11), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT70), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n292), .B2(G68), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT12), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n240), .B1(new_n249), .B2(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n294), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT69), .ZN(new_n416));
  OAI21_X1  g0216(.A(G226), .B1(new_n317), .B2(new_n318), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n268), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n262), .A2(new_n316), .A3(KEYINPUT69), .A4(G226), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n315), .A2(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n271), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n252), .B1(new_n321), .B2(new_n255), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n415), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g0226(.A(KEYINPUT13), .B(new_n424), .C1(new_n422), .C2(new_n271), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n414), .B1(new_n428), .B2(G190), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT71), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n423), .A2(new_n415), .A3(new_n425), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(G190), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n431), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT14), .B1(new_n428), .B2(new_n303), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(G179), .A3(new_n435), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(G169), .C1(new_n426), .C2(new_n427), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n414), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n336), .A2(new_n402), .A3(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n322), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT79), .ZN(new_n450));
  OAI21_X1  g0250(.A(G244), .B1(new_n317), .B2(new_n318), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT4), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G244), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n260), .B2(new_n261), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n316), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n451), .B2(new_n268), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n449), .A2(new_n453), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n271), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n249), .B(G45), .C1(new_n462), .C2(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT80), .B1(new_n462), .B2(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n248), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(G41), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n471), .A2(new_n467), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n254), .A2(G274), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT81), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n271), .B1(new_n465), .B2(new_n467), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n468), .A2(new_n477), .B1(new_n478), .B2(G257), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n460), .A2(new_n461), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(G169), .B1(new_n460), .B2(new_n479), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n293), .A2(new_n206), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n249), .A2(G33), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n292), .A2(new_n483), .A3(new_n278), .A4(new_n277), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n484), .B2(new_n206), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n337), .B2(new_n339), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n285), .A2(KEYINPUT77), .A3(G77), .ZN(new_n487));
  XOR2_X1   g0287(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n488));
  NAND2_X1  g0288(.A1(new_n207), .A2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n208), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(G20), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n286), .B2(new_n204), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n486), .A2(new_n487), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n485), .B1(new_n497), .B2(new_n279), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n480), .A2(new_n481), .A3(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n460), .A2(new_n274), .A3(new_n479), .ZN(new_n500));
  AOI21_X1  g0300(.A(G200), .B1(new_n460), .B2(new_n479), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT82), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n249), .A2(G45), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G250), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n271), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT83), .B1(new_n476), .B2(new_n507), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n248), .A2(new_n511), .A3(new_n473), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n265), .A2(new_n267), .A3(G238), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G244), .A2(G1698), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n319), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n271), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n303), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n519), .A3(new_n461), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n280), .B1(new_n421), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G87), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n206), .A3(new_n207), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n280), .B(G68), .C1(new_n317), .C2(new_n318), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n523), .B1(new_n289), .B2(new_n206), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n279), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n309), .A2(new_n293), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n309), .C2(new_n484), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n521), .A2(new_n522), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n514), .A2(new_n515), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n262), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n254), .B1(new_n536), .B2(new_n517), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n511), .B1(new_n248), .B2(new_n473), .ZN(new_n538));
  AND4_X1   g0338(.A1(new_n511), .A2(new_n254), .A3(G274), .A4(new_n473), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n271), .B2(new_n508), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n513), .A2(new_n519), .A3(G190), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n484), .A2(new_n525), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n531), .A2(new_n532), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n506), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n293), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n313), .A2(G116), .A3(new_n292), .A4(new_n483), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n277), .A2(new_n278), .B1(G20), .B2(new_n549), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(G33), .B2(G283), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G33), .B2(new_n206), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT20), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n262), .A2(new_n316), .A3(G257), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT85), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n322), .A2(G264), .B1(new_n319), .B2(G303), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n254), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n477), .A2(new_n468), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n478), .A2(G270), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT84), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT84), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n388), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n557), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G200), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n568), .ZN(new_n572));
  OR3_X1    g0372(.A1(new_n292), .A2(KEYINPUT25), .A3(G107), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT25), .B1(new_n292), .B2(G107), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n207), .C2(new_n484), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT86), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n280), .B2(G107), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(new_n518), .B2(new_n280), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n262), .A2(new_n280), .A3(G87), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n585), .A2(KEYINPUT24), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n279), .B1(new_n585), .B2(KEYINPUT24), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n576), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n316), .A2(G250), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G257), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n319), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G294), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n259), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n590), .B(new_n271), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n475), .A2(G264), .A3(new_n254), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n562), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n316), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n599), .A2(new_n319), .B1(new_n259), .B2(new_n594), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n590), .B1(new_n600), .B2(new_n271), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n589), .B(G169), .C1(new_n598), .C2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n562), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n271), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(G179), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(KEYINPUT87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n603), .A3(new_n596), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n589), .B1(new_n608), .B2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n588), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n550), .B1(new_n484), .B2(new_n549), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n552), .A2(new_n554), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT20), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(KEYINPUT21), .A3(new_n303), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n557), .B2(G169), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n558), .B(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n560), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n271), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT84), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT84), .B1(new_n562), .B2(new_n563), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT21), .B1(new_n616), .B2(new_n461), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n629), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n604), .A2(new_n562), .A3(new_n597), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n571), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n608), .B2(G190), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n576), .C1(new_n586), .C2(new_n587), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n572), .A2(new_n610), .A3(new_n632), .A4(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n448), .A2(new_n548), .A3(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n448), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT21), .B1(new_n616), .B2(new_n303), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n557), .A2(new_n618), .A3(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n630), .C1(new_n568), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n628), .B2(new_n630), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n610), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(new_n506), .A3(new_n547), .A4(new_n636), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT26), .B1(new_n547), .B2(new_n499), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n460), .A2(new_n479), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n303), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n497), .A2(new_n279), .ZN(new_n652));
  INV_X1    g0452(.A(new_n485), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n460), .A2(new_n461), .A3(new_n479), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n546), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n534), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT90), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT90), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n534), .C1(new_n649), .C2(new_n658), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n648), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n639), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT91), .ZN(new_n665));
  INV_X1    g0465(.A(new_n446), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n440), .B2(new_n331), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT17), .B1(new_n397), .B2(new_n393), .ZN(new_n668));
  INV_X1    g0468(.A(new_n400), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n387), .A2(new_n399), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n302), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n665), .A2(new_n305), .A3(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n249), .A2(new_n280), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n588), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT92), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n610), .A2(new_n636), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n680), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n610), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n616), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n572), .A2(new_n632), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n645), .A2(new_n646), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n632), .A2(new_n680), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n682), .A2(new_n683), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n610), .A2(new_n680), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0501(.A(new_n211), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n526), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n216), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n708));
  XNOR2_X1  g0508(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n663), .A2(new_n685), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n610), .A2(new_n632), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n506), .A3(new_n547), .A4(new_n636), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n534), .B(KEYINPUT96), .Z(new_n714));
  OAI21_X1  g0514(.A(new_n657), .B1(new_n656), .B2(new_n546), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n547), .A2(new_n499), .A3(KEYINPUT26), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n685), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G250), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n592), .B1(new_n268), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n595), .B1(new_n723), .B2(new_n262), .ZN(new_n724));
  OAI211_X1 g0524(.A(G179), .B(new_n597), .C1(new_n724), .C2(new_n254), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(new_n520), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n627), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n460), .A2(new_n479), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT30), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n725), .A2(new_n520), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n730), .B(new_n624), .C1(new_n626), .C2(new_n625), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n650), .A2(new_n461), .A3(new_n633), .A4(new_n520), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n731), .A2(new_n732), .B1(new_n733), .B2(new_n568), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n680), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT31), .B(new_n680), .C1(new_n729), .C2(new_n734), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n506), .A2(new_n547), .A3(new_n685), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n637), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(KEYINPUT95), .A3(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n721), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n709), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n694), .ZN(new_n748));
  INV_X1    g0548(.A(G13), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n249), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n703), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n693), .ZN(new_n755));
  INV_X1    g0555(.A(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n702), .A2(new_n319), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT97), .ZN(new_n758));
  XOR2_X1   g0558(.A(G355), .B(KEYINPUT98), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n244), .A2(new_n472), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n702), .A2(new_n262), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G45), .B2(new_n216), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n760), .B1(G116), .B2(new_n211), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n278), .B1(G20), .B2(new_n303), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n756), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT99), .ZN(new_n771));
  INV_X1    g0571(.A(new_n768), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n461), .A2(new_n571), .A3(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n280), .A2(new_n274), .A3(new_n571), .A4(G179), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n262), .B1(new_n775), .B2(new_n206), .C1(new_n777), .C2(new_n525), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n274), .A2(G20), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT102), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n781), .A2(G179), .A3(new_n571), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n207), .ZN(new_n784));
  NAND2_X1  g0584(.A1(G20), .A2(G179), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT100), .Z(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G200), .A3(new_n569), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n778), .B(new_n784), .C1(G50), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n786), .A2(new_n571), .A3(new_n569), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT101), .Z(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G58), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n786), .A2(new_n274), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n571), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(G200), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G68), .A2(new_n795), .B1(new_n796), .B2(G77), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n781), .A2(G179), .A3(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G159), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT32), .Z(new_n800));
  NAND4_X1  g0600(.A1(new_n789), .A2(new_n793), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  INV_X1    g0602(.A(G326), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n783), .A2(new_n802), .B1(new_n803), .B2(new_n787), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G329), .B2(new_n798), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(G311), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n319), .B1(new_n775), .B2(new_n594), .C1(new_n777), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n790), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G322), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n805), .A2(new_n807), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n772), .B1(new_n801), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n770), .A2(KEYINPUT99), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n767), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n771), .B(new_n816), .C1(new_n693), .C2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n755), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n331), .A2(new_n685), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n333), .A2(new_n334), .B1(new_n314), .B2(new_n680), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n331), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n766), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n594), .A2(new_n790), .B1(new_n787), .B2(new_n809), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n319), .B1(new_n775), .B2(new_n206), .C1(new_n777), .C2(new_n207), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G87), .B2(new_n782), .ZN(new_n828));
  INV_X1    g0628(.A(new_n796), .ZN(new_n829));
  INV_X1    g0629(.A(new_n795), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n549), .B2(new_n829), .C1(new_n802), .C2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n826), .B(new_n831), .C1(G311), .C2(new_n798), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n795), .A2(G150), .B1(new_n788), .B2(G137), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n341), .B2(new_n829), .C1(new_n791), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n262), .B1(new_n777), .B2(new_n238), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G58), .B2(new_n774), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  INV_X1    g0639(.A(new_n798), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n240), .B2(new_n783), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT103), .Z(new_n842));
  AOI21_X1  g0642(.A(new_n832), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n768), .A2(new_n765), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n843), .A2(new_n772), .B1(G77), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n753), .B1(new_n825), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n710), .A2(new_n823), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n663), .A2(new_n685), .A3(new_n824), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(new_n745), .Z(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n851), .B2(new_n753), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(KEYINPUT104), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(KEYINPUT104), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  NOR2_X1   g0656(.A1(new_n750), .A2(new_n249), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n448), .B1(new_n711), .B2(new_n720), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n673), .A2(new_n305), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT107), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n821), .B(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n849), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  INV_X1    g0664(.A(new_n352), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n340), .A2(new_n350), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n345), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n351), .A2(new_n279), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n367), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n678), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n669), .A2(new_n668), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n671), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n386), .B2(new_n870), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n394), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n363), .A2(new_n367), .A3(new_n393), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n363), .A2(new_n367), .B1(new_n384), .B2(new_n385), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n678), .B1(new_n363), .B2(new_n367), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n876), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n864), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n871), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n401), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n368), .A2(new_n386), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n368), .A2(new_n870), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n874), .A4(new_n394), .ZN(new_n887));
  INV_X1    g0687(.A(new_n876), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n414), .A2(new_n680), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n440), .A2(new_n446), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n863), .A2(new_n891), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n879), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n887), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n401), .A2(new_n879), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n903), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n666), .A2(new_n685), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n672), .A2(new_n678), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n902), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n861), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(G330), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n639), .A2(new_n740), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT109), .Z(new_n921));
  NAND4_X1  g0721(.A1(new_n901), .A2(new_n740), .A3(KEYINPUT40), .A4(new_n824), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n909), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n890), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT108), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n904), .A2(new_n909), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n823), .B1(new_n898), .B2(new_n900), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n884), .B2(new_n889), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n740), .B(new_n931), .C1(new_n904), .C2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n926), .A2(new_n929), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n919), .B1(new_n921), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n921), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n857), .B1(new_n918), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n918), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n215), .A2(new_n549), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n490), .A2(new_n493), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT35), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT36), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n343), .A2(G77), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n239), .B1(new_n216), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n749), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n944), .A3(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n654), .A2(new_n680), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n506), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT110), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n499), .A2(new_n680), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n954), .A2(new_n683), .A3(new_n682), .A4(new_n696), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n656), .B1(new_n952), .B2(new_n610), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n955), .A2(KEYINPUT42), .B1(new_n957), .B2(new_n685), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n544), .A2(new_n685), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n547), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n534), .A2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n695), .A2(new_n954), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n956), .A2(new_n958), .A3(new_n965), .A4(new_n964), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n703), .B(new_n974), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n695), .ZN(new_n977));
  AND2_X1   g0777(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n952), .A2(new_n699), .A3(new_n953), .ZN(new_n979));
  NOR2_X1   g0779(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n699), .B1(new_n952), .B2(new_n953), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT45), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n977), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n697), .B1(new_n687), .B2(new_n696), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n748), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n721), .A2(new_n745), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n982), .A2(new_n984), .A3(new_n977), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n976), .B1(new_n991), .B2(new_n746), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n973), .B1(new_n992), .B2(new_n752), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n233), .A2(new_n762), .ZN(new_n994));
  INV_X1    g0794(.A(new_n309), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n768), .B(new_n767), .C1(new_n702), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n756), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT115), .B(G137), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n798), .A2(new_n999), .B1(G58), .B2(new_n776), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT116), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n782), .A2(G77), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n262), .C1(new_n834), .C2(new_n787), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n238), .A2(new_n829), .B1(new_n830), .B2(new_n341), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n790), .A2(new_n287), .B1(new_n240), .B2(new_n775), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT114), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n776), .A2(G116), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1008), .A2(new_n1009), .B1(G107), .B2(new_n774), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G311), .B2(new_n788), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G283), .A2(new_n796), .B1(new_n795), .B2(G294), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n809), .C2(new_n791), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n782), .A2(G97), .ZN(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n319), .C1(new_n840), .C2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT113), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1005), .A2(new_n1007), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n997), .B1(new_n817), .B2(new_n963), .C1(new_n1020), .C2(new_n772), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n993), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n752), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n230), .A2(new_n472), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n705), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1024), .A2(new_n762), .B1(new_n1025), .B2(new_n758), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n705), .B(new_n472), .C1(new_n240), .C2(new_n204), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n311), .B2(new_n238), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n288), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1026), .A2(new_n1031), .B1(G107), .B2(new_n211), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n756), .B1(new_n1032), .B2(new_n769), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n777), .A2(new_n204), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n319), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1015), .B(new_n1035), .C1(new_n840), .C2(new_n287), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT117), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n995), .A2(new_n774), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n787), .B2(new_n341), .C1(new_n238), .C2(new_n790), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n240), .A2(new_n829), .B1(new_n830), .B2(new_n288), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n795), .A2(G311), .B1(new_n788), .B2(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n809), .B2(new_n829), .C1(new_n791), .C2(new_n1016), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n776), .A2(G294), .B1(new_n774), .B2(G283), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n319), .B1(new_n783), .B2(new_n549), .C1(new_n803), .C2(new_n840), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1049), .B2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1041), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1033), .B1(new_n687), .B2(new_n817), .C1(new_n1053), .C2(new_n772), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n989), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n703), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n746), .A2(new_n988), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1023), .B(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  INV_X1    g0858(.A(new_n990), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1059), .A2(new_n751), .A3(new_n985), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n952), .A2(new_n767), .A3(new_n953), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n762), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n769), .B1(new_n206), .B2(new_n211), .C1(new_n237), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n753), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n811), .B1(new_n788), .B2(G317), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT52), .Z(new_n1066));
  OAI221_X1 g0866(.A(new_n319), .B1(new_n775), .B2(new_n549), .C1(new_n777), .C2(new_n802), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1067), .B(new_n784), .C1(G322), .C2(new_n798), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G294), .A2(new_n796), .B1(new_n795), .B2(G303), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n796), .A2(new_n311), .B1(G77), .B2(new_n774), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n238), .B2(new_n830), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT118), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n287), .A2(new_n787), .B1(new_n790), .B2(new_n341), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n782), .A2(G87), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n798), .A2(G143), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n319), .B1(new_n776), .B2(G68), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1070), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1064), .B1(new_n1080), .B2(new_n768), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1060), .B1(new_n1061), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1055), .B1(new_n1059), .B2(new_n985), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n703), .A3(new_n991), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(G390));
  NAND2_X1  g0885(.A1(new_n910), .A2(new_n911), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n898), .A2(new_n900), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n849), .B2(new_n862), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1088), .B2(new_n913), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n718), .A2(new_n824), .A3(new_n685), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1087), .B1(new_n1090), .B2(new_n862), .ZN(new_n1091));
  OR3_X1    g0891(.A1(new_n1091), .A2(new_n928), .A3(new_n913), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n743), .A2(new_n744), .A3(new_n824), .A4(new_n901), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1091), .A2(new_n928), .A3(new_n913), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n863), .A2(new_n901), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n912), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1095), .B1(new_n1097), .B2(new_n1086), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n741), .A2(new_n1087), .A3(new_n823), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1094), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1090), .A2(new_n862), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n740), .A2(G330), .A3(new_n824), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1087), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1093), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n743), .A2(new_n744), .A3(new_n824), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1099), .B1(new_n1106), .B2(new_n1087), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n863), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n448), .A2(new_n741), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n858), .A2(new_n859), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1096), .A2(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1099), .B1(new_n1114), .B2(new_n1095), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1115), .A2(new_n1109), .A3(new_n1111), .A4(new_n1094), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n703), .A3(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1115), .A2(new_n1094), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1086), .A2(new_n765), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n753), .B1(new_n311), .B2(new_n845), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n840), .A2(new_n594), .B1(new_n802), .B2(new_n787), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n262), .B1(new_n776), .B2(G87), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(KEYINPUT121), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n782), .A2(G68), .B1(G77), .B2(new_n774), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G116), .B2(new_n811), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G97), .A2(new_n796), .B1(new_n795), .B2(G107), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1129), .A2(new_n787), .B1(new_n790), .B2(new_n839), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT120), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n795), .A2(new_n999), .B1(new_n796), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n776), .A2(G150), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1137), .A2(KEYINPUT53), .B1(new_n341), .B2(new_n775), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n319), .B(new_n1138), .C1(KEYINPUT53), .C2(new_n1137), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G50), .A2(new_n782), .B1(new_n798), .B2(G125), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(KEYINPUT119), .C2(new_n1134), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1128), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1120), .B1(new_n1142), .B2(new_n768), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1118), .A2(new_n752), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1117), .B1(new_n1145), .B2(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT125), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n297), .A2(new_n870), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n306), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1150), .B(new_n1151), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n919), .B1(new_n933), .B2(new_n930), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT108), .B1(new_n923), .B2(new_n925), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n928), .A2(new_n922), .A3(new_n927), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n917), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n926), .A2(new_n929), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n916), .B1(new_n1159), .B2(new_n1154), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1153), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n917), .A2(new_n1157), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n916), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1152), .A3(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1161), .A2(new_n1164), .B1(new_n1116), .B2(new_n1111), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1148), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n704), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1109), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1111), .B1(new_n1101), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1164), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(KEYINPUT125), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1166), .A2(new_n1167), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n751), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n765), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n753), .B1(G50), .B2(new_n845), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G132), .A2(new_n795), .B1(new_n796), .B2(G137), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT123), .Z(new_n1180));
  AOI22_X1  g0980(.A1(G125), .A2(new_n788), .B1(new_n811), .B2(G128), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n776), .A2(new_n1133), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT124), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n287), .C2(new_n775), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n259), .B(new_n462), .C1(new_n783), .C2(new_n341), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G124), .B2(new_n798), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n788), .A2(G116), .B1(new_n782), .B2(G58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n207), .B2(new_n790), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n319), .A2(new_n462), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1034), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n240), .B2(new_n775), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G283), .B2(new_n798), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n206), .B2(new_n830), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1193), .B(new_n1198), .C1(new_n995), .C2(new_n796), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1194), .B(new_n238), .C1(G33), .C2(G41), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1191), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1178), .B1(new_n1203), .B2(new_n768), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1176), .B1(new_n1177), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1175), .A2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1109), .A2(new_n752), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n287), .A2(new_n829), .B1(new_n830), .B2(new_n1132), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n262), .B1(new_n775), .B2(new_n238), .C1(new_n777), .C2(new_n341), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G58), .B2(new_n782), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n1129), .B2(new_n840), .C1(new_n839), .C2(new_n787), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(new_n792), .C2(new_n999), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n795), .A2(G116), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n262), .B1(new_n776), .B2(G97), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n1002), .A3(new_n1038), .A4(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G283), .A2(new_n811), .B1(new_n788), .B2(G294), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n809), .B2(new_n840), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G107), .C2(new_n796), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n768), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n756), .B1(new_n240), .B2(new_n844), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n901), .C2(new_n766), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1207), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT126), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n975), .A3(new_n1112), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(G381));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1227), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1144), .A2(new_n1117), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G375), .A2(new_n1228), .A3(G381), .A4(new_n1230), .ZN(G407));
  NAND2_X1  g1031(.A1(new_n679), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G375), .C2(new_n1234), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1175), .A2(G378), .A3(new_n1205), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1205), .B1(new_n976), .B2(new_n1172), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1229), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1109), .A2(new_n1111), .A3(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(new_n704), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1224), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n855), .B1(new_n1223), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1223), .A2(new_n1246), .A3(new_n855), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1233), .A2(G2897), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1249), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1253), .B2(new_n1247), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1236), .B1(new_n1240), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1232), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1253), .A2(new_n1247), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(new_n819), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n993), .B2(new_n1021), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n993), .A2(G390), .A3(new_n1021), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1264), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(KEYINPUT127), .B(new_n1263), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1261), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1257), .A2(new_n1262), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1240), .A2(new_n1276), .A3(new_n1273), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1240), .B2(new_n1273), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1277), .A2(new_n1256), .A3(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1279), .B2(new_n1272), .ZN(G405));
  OAI21_X1  g1080(.A(new_n1261), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1229), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(new_n1237), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1268), .A2(new_n1269), .A3(new_n1264), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1267), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1269), .B1(new_n1285), .B2(new_n1265), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1263), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1287), .A3(new_n1273), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1281), .A2(new_n1283), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1283), .B1(new_n1281), .B2(new_n1288), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(G402));
endmodule


