

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718;

  AND2_X1 U372 ( .A1(n711), .A2(n412), .ZN(n411) );
  XNOR2_X1 U373 ( .A(n471), .B(n423), .ZN(n491) );
  NAND2_X1 U374 ( .A1(n421), .A2(n422), .ZN(n389) );
  INV_X1 U375 ( .A(G143), .ZN(n419) );
  INV_X2 U376 ( .A(G953), .ZN(n705) );
  XNOR2_X2 U377 ( .A(n698), .B(n505), .ZN(n676) );
  NAND2_X2 U378 ( .A1(n408), .A2(n360), .ZN(n409) );
  XNOR2_X1 U379 ( .A(KEYINPUT72), .B(G119), .ZN(n370) );
  XNOR2_X1 U380 ( .A(G104), .B(G110), .ZN(n483) );
  XNOR2_X1 U381 ( .A(n407), .B(n406), .ZN(n578) );
  XNOR2_X1 U382 ( .A(n572), .B(KEYINPUT32), .ZN(n364) );
  XNOR2_X1 U383 ( .A(KEYINPUT106), .B(n570), .ZN(n712) );
  AND2_X4 U384 ( .A1(n409), .A2(n595), .ZN(n681) );
  XNOR2_X2 U385 ( .A(n504), .B(n503), .ZN(n698) );
  XNOR2_X2 U386 ( .A(n496), .B(n495), .ZN(n545) );
  INV_X1 U387 ( .A(n645), .ZN(n576) );
  XNOR2_X1 U388 ( .A(n387), .B(n410), .ZN(n386) );
  NOR2_X1 U389 ( .A1(n648), .A2(n647), .ZN(n372) );
  NOR2_X1 U390 ( .A1(n363), .A2(n647), .ZN(n581) );
  XNOR2_X1 U391 ( .A(n453), .B(n452), .ZN(n645) );
  XNOR2_X2 U392 ( .A(KEYINPUT10), .B(n443), .ZN(n697) );
  NAND2_X1 U393 ( .A1(n386), .A2(n418), .ZN(n385) );
  AND2_X2 U394 ( .A1(n712), .A2(n364), .ZN(n588) );
  NOR2_X1 U395 ( .A1(n390), .A2(n559), .ZN(n560) );
  INV_X1 U396 ( .A(n567), .ZN(n352) );
  XNOR2_X1 U397 ( .A(n372), .B(KEYINPUT75), .ZN(n577) );
  INV_X1 U398 ( .A(n509), .ZN(n510) );
  XNOR2_X1 U399 ( .A(G116), .B(G101), .ZN(n430) );
  XNOR2_X1 U400 ( .A(G113), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X1 U401 ( .A(n362), .B(KEYINPUT33), .ZN(n390) );
  NOR2_X1 U402 ( .A1(n577), .A2(n353), .ZN(n362) );
  XNOR2_X1 U403 ( .A(n518), .B(n507), .ZN(n648) );
  XNOR2_X1 U404 ( .A(n506), .B(G469), .ZN(n518) );
  XNOR2_X1 U405 ( .A(n369), .B(n368), .ZN(n486) );
  XNOR2_X1 U406 ( .A(n430), .B(n370), .ZN(n369) );
  XNOR2_X1 U407 ( .A(n431), .B(KEYINPUT71), .ZN(n368) );
  NOR2_X1 U408 ( .A1(n676), .A2(G902), .ZN(n506) );
  XNOR2_X1 U409 ( .A(n486), .B(n485), .ZN(n686) );
  XNOR2_X1 U410 ( .A(n502), .B(n484), .ZN(n485) );
  XOR2_X1 U411 ( .A(G122), .B(KEYINPUT16), .Z(n484) );
  NAND2_X1 U412 ( .A1(n545), .A2(n635), .ZN(n521) );
  XNOR2_X1 U413 ( .A(n491), .B(n425), .ZN(n504) );
  XNOR2_X1 U414 ( .A(n424), .B(G134), .ZN(n425) );
  XOR2_X1 U415 ( .A(KEYINPUT70), .B(G131), .Z(n424) );
  XOR2_X1 U416 ( .A(G137), .B(G140), .Z(n503) );
  XNOR2_X1 U417 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U418 ( .A1(n670), .A2(n590), .ZN(n496) );
  XOR2_X1 U419 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n459) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT100), .ZN(n458) );
  XOR2_X1 U421 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n457) );
  INV_X1 U422 ( .A(KEYINPUT44), .ZN(n412) );
  OR2_X1 U423 ( .A1(G237), .A2(G902), .ZN(n497) );
  NOR2_X1 U424 ( .A1(n454), .A2(n513), .ZN(n517) );
  NOR2_X1 U425 ( .A1(n634), .A2(n566), .ZN(n405) );
  XNOR2_X1 U426 ( .A(n361), .B(n504), .ZN(n480) );
  XNOR2_X1 U427 ( .A(n434), .B(n429), .ZN(n361) );
  XNOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n379) );
  XNOR2_X1 U429 ( .A(G119), .B(G128), .ZN(n444) );
  XOR2_X1 U430 ( .A(KEYINPUT23), .B(G110), .Z(n445) );
  XOR2_X1 U431 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n469) );
  XNOR2_X1 U432 ( .A(G134), .B(KEYINPUT9), .ZN(n468) );
  XNOR2_X1 U433 ( .A(G116), .B(G107), .ZN(n473) );
  XOR2_X1 U434 ( .A(KEYINPUT101), .B(G122), .Z(n474) );
  XNOR2_X1 U435 ( .A(n465), .B(n400), .ZN(n602) );
  XNOR2_X1 U436 ( .A(n697), .B(n401), .ZN(n400) );
  XNOR2_X1 U437 ( .A(n455), .B(n402), .ZN(n401) );
  INV_X1 U438 ( .A(KEYINPUT0), .ZN(n406) );
  NAND2_X1 U439 ( .A1(n558), .A2(n557), .ZN(n407) );
  XNOR2_X1 U440 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U441 ( .A1(G902), .A2(n683), .ZN(n453) );
  XNOR2_X1 U442 ( .A(n416), .B(n414), .ZN(n490) );
  XNOR2_X1 U443 ( .A(n489), .B(n415), .ZN(n414) );
  NOR2_X1 U444 ( .A1(G952), .A2(n705), .ZN(n685) );
  XNOR2_X1 U445 ( .A(n630), .B(KEYINPUT84), .ZN(n631) );
  NOR2_X1 U446 ( .A1(n354), .A2(n371), .ZN(n393) );
  NOR2_X1 U447 ( .A1(KEYINPUT69), .A2(n525), .ZN(n526) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n432) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U450 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n426) );
  XOR2_X1 U451 ( .A(G146), .B(G137), .Z(n427) );
  INV_X1 U452 ( .A(G128), .ZN(n420) );
  XNOR2_X1 U453 ( .A(G113), .B(G131), .ZN(n455) );
  INV_X1 U454 ( .A(G104), .ZN(n402) );
  XNOR2_X1 U455 ( .A(G143), .B(G122), .ZN(n456) );
  XNOR2_X1 U456 ( .A(n588), .B(n587), .ZN(n413) );
  INV_X1 U457 ( .A(KEYINPUT87), .ZN(n587) );
  INV_X1 U458 ( .A(KEYINPUT73), .ZN(n410) );
  NAND2_X1 U459 ( .A1(G234), .A2(G237), .ZN(n435) );
  NAND2_X1 U460 ( .A1(n517), .A2(n654), .ZN(n384) );
  XNOR2_X1 U461 ( .A(n521), .B(n520), .ZN(n558) );
  BUF_X1 U462 ( .A(n518), .Z(n363) );
  XOR2_X1 U463 ( .A(G101), .B(G146), .Z(n500) );
  INV_X1 U464 ( .A(KEYINPUT4), .ZN(n423) );
  XNOR2_X1 U465 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n415) );
  XNOR2_X1 U466 ( .A(n488), .B(n487), .ZN(n416) );
  INV_X1 U467 ( .A(KEYINPUT86), .ZN(n551) );
  AND2_X1 U468 ( .A1(n382), .A2(n381), .ZN(n535) );
  INV_X1 U469 ( .A(n363), .ZN(n381) );
  XNOR2_X1 U470 ( .A(n384), .B(n383), .ZN(n382) );
  INV_X1 U471 ( .A(KEYINPUT28), .ZN(n383) );
  INV_X1 U472 ( .A(n635), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n530), .B(n529), .ZN(n548) );
  NOR2_X1 U474 ( .A1(n528), .A2(n632), .ZN(n530) );
  XNOR2_X1 U475 ( .A(n403), .B(n367), .ZN(n366) );
  INV_X1 U476 ( .A(KEYINPUT22), .ZN(n367) );
  XNOR2_X1 U477 ( .A(n405), .B(KEYINPUT104), .ZN(n404) );
  NOR2_X1 U478 ( .A1(n602), .A2(G902), .ZN(n467) );
  AND2_X1 U479 ( .A1(n366), .A2(n353), .ZN(n574) );
  XNOR2_X1 U480 ( .A(n596), .B(n597), .ZN(n598) );
  XNOR2_X1 U481 ( .A(n448), .B(n377), .ZN(n683) );
  XNOR2_X1 U482 ( .A(n380), .B(n378), .ZN(n377) );
  XNOR2_X1 U483 ( .A(n503), .B(n379), .ZN(n378) );
  XNOR2_X1 U484 ( .A(n476), .B(n477), .ZN(n679) );
  XNOR2_X1 U485 ( .A(n602), .B(KEYINPUT59), .ZN(n603) );
  NAND2_X1 U486 ( .A1(n681), .A2(G475), .ZN(n604) );
  NOR2_X1 U487 ( .A1(n542), .A2(n521), .ZN(n498) );
  NOR2_X1 U488 ( .A1(n547), .A2(n524), .ZN(n617) );
  NOR2_X1 U489 ( .A1(n533), .A2(n523), .ZN(n622) );
  XNOR2_X1 U490 ( .A(n399), .B(n398), .ZN(n677) );
  XNOR2_X1 U491 ( .A(n676), .B(n675), .ZN(n398) );
  XNOR2_X1 U492 ( .A(n671), .B(n672), .ZN(n673) );
  AND2_X1 U493 ( .A1(n665), .A2(n705), .ZN(n391) );
  NAND2_X1 U494 ( .A1(n631), .A2(n393), .ZN(n392) );
  XNOR2_X1 U495 ( .A(n654), .B(KEYINPUT6), .ZN(n353) );
  NOR2_X1 U496 ( .A1(n703), .A2(KEYINPUT2), .ZN(n354) );
  XOR2_X1 U497 ( .A(KEYINPUT105), .B(n585), .Z(n355) );
  AND2_X1 U498 ( .A1(n629), .A2(n620), .ZN(n356) );
  NOR2_X1 U499 ( .A1(n642), .A2(n390), .ZN(n357) );
  AND2_X1 U500 ( .A1(n550), .A2(n716), .ZN(n358) );
  NOR2_X1 U501 ( .A1(n390), .A2(n663), .ZN(n359) );
  OR2_X1 U502 ( .A1(n592), .A2(n591), .ZN(n360) );
  XOR2_X1 U503 ( .A(G902), .B(KEYINPUT15), .Z(n590) );
  INV_X1 U504 ( .A(n443), .ZN(n488) );
  NOR2_X1 U505 ( .A1(n679), .A2(G902), .ZN(n478) );
  INV_X1 U506 ( .A(n509), .ZN(n654) );
  XNOR2_X1 U507 ( .A(n375), .B(n374), .ZN(n373) );
  NAND2_X1 U508 ( .A1(n373), .A2(n358), .ZN(n593) );
  XNOR2_X1 U509 ( .A(n364), .B(G119), .ZN(n709) );
  NAND2_X1 U510 ( .A1(n589), .A2(n365), .ZN(n408) );
  NAND2_X1 U511 ( .A1(n365), .A2(n594), .ZN(n595) );
  OR2_X1 U512 ( .A1(n365), .A2(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U513 ( .A1(n365), .A2(n705), .ZN(n693) );
  XNOR2_X2 U514 ( .A(n385), .B(KEYINPUT45), .ZN(n365) );
  AND2_X1 U515 ( .A1(n366), .A2(n352), .ZN(n569) );
  INV_X1 U516 ( .A(n595), .ZN(n371) );
  NAND2_X1 U517 ( .A1(n376), .A2(n539), .ZN(n375) );
  AND2_X1 U518 ( .A1(n356), .A2(n540), .ZN(n376) );
  NAND2_X1 U519 ( .A1(n472), .A2(G221), .ZN(n380) );
  NAND2_X1 U520 ( .A1(n411), .A2(n413), .ZN(n387) );
  XNOR2_X2 U521 ( .A(n389), .B(n388), .ZN(n471) );
  XNOR2_X2 U522 ( .A(KEYINPUT65), .B(KEYINPUT81), .ZN(n388) );
  NAND2_X1 U523 ( .A1(n392), .A2(n391), .ZN(n666) );
  XNOR2_X2 U524 ( .A(G146), .B(G125), .ZN(n443) );
  XNOR2_X1 U525 ( .A(n394), .B(KEYINPUT41), .ZN(n643) );
  NAND2_X1 U526 ( .A1(n397), .A2(n395), .ZN(n394) );
  NOR2_X1 U527 ( .A1(n634), .A2(n396), .ZN(n395) );
  INV_X1 U528 ( .A(n632), .ZN(n397) );
  NAND2_X1 U529 ( .A1(n681), .A2(G469), .ZN(n399) );
  NAND2_X1 U530 ( .A1(n578), .A2(n404), .ZN(n403) );
  XNOR2_X1 U531 ( .A(n490), .B(n491), .ZN(n492) );
  XOR2_X1 U532 ( .A(n474), .B(n473), .Z(n417) );
  AND2_X1 U533 ( .A1(n586), .A2(n355), .ZN(n418) );
  XNOR2_X1 U534 ( .A(n428), .B(KEYINPUT76), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n486), .B(n433), .ZN(n434) );
  XNOR2_X1 U536 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U537 ( .A(KEYINPUT39), .ZN(n529) );
  INV_X1 U538 ( .A(KEYINPUT91), .ZN(n493) );
  XNOR2_X1 U539 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U540 ( .A(n599), .B(KEYINPUT63), .ZN(n600) );
  XNOR2_X1 U541 ( .A(KEYINPUT60), .B(KEYINPUT68), .ZN(n607) );
  XNOR2_X1 U542 ( .A(n532), .B(n531), .ZN(n715) );
  NAND2_X1 U543 ( .A1(n419), .A2(G128), .ZN(n422) );
  NAND2_X1 U544 ( .A1(n420), .A2(G143), .ZN(n421) );
  XNOR2_X1 U545 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U546 ( .A(KEYINPUT77), .B(n432), .Z(n462) );
  NAND2_X1 U547 ( .A1(n462), .A2(G210), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n480), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U549 ( .A(n435), .B(KEYINPUT14), .ZN(n436) );
  NAND2_X1 U550 ( .A1(G952), .A2(n436), .ZN(n662) );
  NOR2_X1 U551 ( .A1(G953), .A2(n662), .ZN(n556) );
  NAND2_X1 U552 ( .A1(n436), .A2(G902), .ZN(n437) );
  XOR2_X1 U553 ( .A(KEYINPUT92), .B(n437), .Z(n553) );
  NAND2_X1 U554 ( .A1(n553), .A2(G953), .ZN(n438) );
  NOR2_X1 U555 ( .A1(G900), .A2(n438), .ZN(n439) );
  NOR2_X1 U556 ( .A1(n556), .A2(n439), .ZN(n513) );
  INV_X1 U557 ( .A(n590), .ZN(n552) );
  NAND2_X1 U558 ( .A1(G234), .A2(n552), .ZN(n440) );
  XNOR2_X1 U559 ( .A(KEYINPUT20), .B(n440), .ZN(n449) );
  NAND2_X1 U560 ( .A1(G221), .A2(n449), .ZN(n441) );
  XOR2_X1 U561 ( .A(KEYINPUT21), .B(n441), .Z(n644) );
  NAND2_X1 U562 ( .A1(G234), .A2(n705), .ZN(n442) );
  XOR2_X1 U563 ( .A(KEYINPUT8), .B(n442), .Z(n472) );
  XNOR2_X1 U564 ( .A(n697), .B(KEYINPUT83), .ZN(n447) );
  XNOR2_X1 U565 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U566 ( .A1(G217), .A2(n449), .ZN(n451) );
  XNOR2_X1 U567 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n450) );
  NAND2_X1 U568 ( .A1(n644), .A2(n576), .ZN(n454) );
  XNOR2_X1 U569 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U571 ( .A(n461), .B(n460), .Z(n464) );
  NAND2_X1 U572 ( .A1(G214), .A2(n462), .ZN(n463) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(G475), .ZN(n466) );
  XOR2_X1 U574 ( .A(n467), .B(n466), .Z(n533) );
  XNOR2_X1 U575 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U576 ( .A(n471), .B(n470), .Z(n477) );
  NAND2_X1 U577 ( .A1(G217), .A2(n472), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n475), .B(n417), .ZN(n476) );
  XOR2_X1 U579 ( .A(G478), .B(n478), .Z(n479) );
  XNOR2_X1 U580 ( .A(n479), .B(KEYINPUT103), .ZN(n534) );
  INV_X1 U581 ( .A(n534), .ZN(n523) );
  INV_X1 U582 ( .A(n622), .ZN(n522) );
  NOR2_X1 U583 ( .A1(G902), .A2(n480), .ZN(n481) );
  XNOR2_X1 U584 ( .A(G472), .B(n481), .ZN(n509) );
  NOR2_X1 U585 ( .A1(n522), .A2(n353), .ZN(n482) );
  NAND2_X1 U586 ( .A1(n517), .A2(n482), .ZN(n542) );
  XNOR2_X1 U587 ( .A(n483), .B(G107), .ZN(n502) );
  XNOR2_X1 U588 ( .A(KEYINPUT90), .B(KEYINPUT79), .ZN(n487) );
  NAND2_X1 U589 ( .A1(G224), .A2(n705), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n686), .B(n492), .ZN(n670) );
  NAND2_X1 U591 ( .A1(G210), .A2(n497), .ZN(n494) );
  NAND2_X1 U592 ( .A1(G214), .A2(n497), .ZN(n635) );
  XNOR2_X1 U593 ( .A(KEYINPUT36), .B(n498), .ZN(n508) );
  XNOR2_X1 U594 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n507) );
  NAND2_X1 U595 ( .A1(G227), .A2(n705), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n505) );
  INV_X1 U598 ( .A(n648), .ZN(n567) );
  NAND2_X1 U599 ( .A1(n508), .A2(n567), .ZN(n629) );
  NAND2_X1 U600 ( .A1(n510), .A2(n635), .ZN(n511) );
  XNOR2_X1 U601 ( .A(n511), .B(KEYINPUT30), .ZN(n512) );
  NOR2_X1 U602 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U603 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U604 ( .A1(n514), .A2(n581), .ZN(n528) );
  OR2_X1 U605 ( .A1(n533), .A2(n534), .ZN(n515) );
  XOR2_X1 U606 ( .A(KEYINPUT107), .B(n515), .Z(n561) );
  NOR2_X1 U607 ( .A1(n528), .A2(n561), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n545), .A2(n516), .ZN(n620) );
  XOR2_X1 U609 ( .A(KEYINPUT78), .B(KEYINPUT19), .Z(n519) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n519), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n535), .A2(n558), .ZN(n524) );
  NOR2_X1 U612 ( .A1(n524), .A2(n522), .ZN(n621) );
  NAND2_X1 U613 ( .A1(n533), .A2(n523), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n621), .A2(n617), .ZN(n525) );
  XNOR2_X1 U615 ( .A(KEYINPUT47), .B(n526), .ZN(n540) );
  XNOR2_X1 U616 ( .A(n545), .B(KEYINPUT38), .ZN(n527) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT74), .ZN(n632) );
  NAND2_X1 U618 ( .A1(n622), .A2(n548), .ZN(n532) );
  XOR2_X1 U619 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n531) );
  NAND2_X1 U620 ( .A1(n534), .A2(n533), .ZN(n634) );
  NAND2_X1 U621 ( .A1(n535), .A2(n643), .ZN(n536) );
  XNOR2_X1 U622 ( .A(n536), .B(KEYINPUT42), .ZN(n717) );
  NAND2_X1 U623 ( .A1(n715), .A2(n717), .ZN(n538) );
  XOR2_X1 U624 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n537) );
  XNOR2_X1 U625 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n635), .A2(n352), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n543), .B(KEYINPUT43), .ZN(n544) );
  NOR2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U630 ( .A(KEYINPUT108), .B(n546), .ZN(n713) );
  INV_X1 U631 ( .A(n713), .ZN(n550) );
  INV_X1 U632 ( .A(n547), .ZN(n624) );
  NAND2_X1 U633 ( .A1(n548), .A2(n624), .ZN(n549) );
  XNOR2_X1 U634 ( .A(KEYINPUT110), .B(n549), .ZN(n716) );
  XNOR2_X2 U635 ( .A(n593), .B(n551), .ZN(n703) );
  AND2_X1 U636 ( .A1(n703), .A2(n590), .ZN(n589) );
  NOR2_X1 U637 ( .A1(G898), .A2(n705), .ZN(n688) );
  NAND2_X1 U638 ( .A1(n688), .A2(n553), .ZN(n554) );
  XNOR2_X1 U639 ( .A(KEYINPUT93), .B(n554), .ZN(n555) );
  OR2_X1 U640 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT94), .ZN(n580) );
  INV_X1 U642 ( .A(n580), .ZN(n559) );
  XNOR2_X1 U643 ( .A(n560), .B(KEYINPUT34), .ZN(n563) );
  XOR2_X1 U644 ( .A(n561), .B(KEYINPUT80), .Z(n562) );
  NAND2_X1 U645 ( .A1(n563), .A2(n562), .ZN(n565) );
  INV_X1 U646 ( .A(KEYINPUT35), .ZN(n564) );
  XNOR2_X2 U647 ( .A(n565), .B(n564), .ZN(n711) );
  INV_X1 U648 ( .A(n644), .ZN(n566) );
  NOR2_X1 U649 ( .A1(n654), .A2(n645), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U651 ( .A1(n352), .A2(n645), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n574), .A2(n571), .ZN(n572) );
  NAND2_X1 U653 ( .A1(n711), .A2(n588), .ZN(n573) );
  NAND2_X1 U654 ( .A1(n573), .A2(KEYINPUT44), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n574), .A2(n352), .ZN(n575) );
  NOR2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n609) );
  NOR2_X1 U657 ( .A1(n624), .A2(n622), .ZN(n637) );
  NOR2_X1 U658 ( .A1(n509), .A2(n577), .ZN(n656) );
  NAND2_X1 U659 ( .A1(n578), .A2(n656), .ZN(n579) );
  XNOR2_X1 U660 ( .A(n579), .B(KEYINPUT31), .ZN(n625) );
  NAND2_X1 U661 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U662 ( .A1(n654), .A2(n582), .ZN(n614) );
  NOR2_X1 U663 ( .A1(n625), .A2(n614), .ZN(n583) );
  NOR2_X1 U664 ( .A1(n637), .A2(n583), .ZN(n584) );
  NOR2_X1 U665 ( .A1(n609), .A2(n584), .ZN(n585) );
  INV_X1 U666 ( .A(KEYINPUT2), .ZN(n592) );
  XNOR2_X1 U667 ( .A(KEYINPUT85), .B(n590), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n681), .A2(G472), .ZN(n596) );
  NOR2_X2 U670 ( .A1(n598), .A2(n685), .ZN(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n601), .B(n600), .ZN(G57) );
  INV_X1 U673 ( .A(n685), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(n605) );
  AND2_X2 U675 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(n607), .ZN(G60) );
  XOR2_X1 U677 ( .A(G101), .B(n609), .Z(G3) );
  NAND2_X1 U678 ( .A1(n614), .A2(n622), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n610), .B(G104), .ZN(G6) );
  XOR2_X1 U680 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n612) );
  XNOR2_X1 U681 ( .A(G107), .B(KEYINPUT26), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT111), .B(n613), .Z(n616) );
  NAND2_X1 U684 ( .A1(n614), .A2(n624), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(G9) );
  XOR2_X1 U686 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n619) );
  XNOR2_X1 U687 ( .A(G128), .B(n617), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(G30) );
  XNOR2_X1 U689 ( .A(G143), .B(n620), .ZN(G45) );
  XOR2_X1 U690 ( .A(G146), .B(n621), .Z(G48) );
  NAND2_X1 U691 ( .A1(n625), .A2(n622), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n623), .B(G113), .ZN(G15) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U694 ( .A(n626), .B(KEYINPUT114), .ZN(n627) );
  XNOR2_X1 U695 ( .A(G116), .B(n627), .ZN(G18) );
  XOR2_X1 U696 ( .A(G125), .B(KEYINPUT37), .Z(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(G27) );
  NOR2_X1 U698 ( .A1(n397), .A2(n635), .ZN(n633) );
  NOR2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n640) );
  NAND2_X1 U700 ( .A1(n397), .A2(n635), .ZN(n636) );
  NOR2_X1 U701 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U702 ( .A(KEYINPUT117), .B(n638), .Z(n639) );
  NOR2_X1 U703 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U704 ( .A(n641), .B(KEYINPUT118), .ZN(n642) );
  INV_X1 U705 ( .A(n643), .ZN(n663) );
  NOR2_X1 U706 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U707 ( .A(KEYINPUT49), .B(n646), .ZN(n652) );
  NAND2_X1 U708 ( .A1(n352), .A2(n647), .ZN(n649) );
  XNOR2_X1 U709 ( .A(n649), .B(KEYINPUT116), .ZN(n650) );
  XNOR2_X1 U710 ( .A(KEYINPUT50), .B(n650), .ZN(n651) );
  NAND2_X1 U711 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U712 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U713 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U714 ( .A(KEYINPUT51), .B(n657), .Z(n658) );
  NOR2_X1 U715 ( .A1(n663), .A2(n658), .ZN(n659) );
  NOR2_X1 U716 ( .A1(n357), .A2(n659), .ZN(n660) );
  XNOR2_X1 U717 ( .A(n660), .B(KEYINPUT52), .ZN(n661) );
  NOR2_X1 U718 ( .A1(n662), .A2(n661), .ZN(n664) );
  NOR2_X1 U719 ( .A1(n664), .A2(n359), .ZN(n665) );
  XOR2_X1 U720 ( .A(KEYINPUT53), .B(n666), .Z(G75) );
  XOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n668) );
  XNOR2_X1 U722 ( .A(KEYINPUT82), .B(KEYINPUT55), .ZN(n667) );
  XNOR2_X1 U723 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U724 ( .A(n670), .B(n669), .Z(n672) );
  NAND2_X1 U725 ( .A1(n681), .A2(G210), .ZN(n671) );
  NOR2_X2 U726 ( .A1(n673), .A2(n685), .ZN(n674) );
  XNOR2_X1 U727 ( .A(n674), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U728 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n675) );
  NOR2_X1 U729 ( .A1(n685), .A2(n677), .ZN(G54) );
  NAND2_X1 U730 ( .A1(G478), .A2(n681), .ZN(n678) );
  XNOR2_X1 U731 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U732 ( .A1(n685), .A2(n680), .ZN(G63) );
  NAND2_X1 U733 ( .A1(G217), .A2(n681), .ZN(n682) );
  XNOR2_X1 U734 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U735 ( .A1(n685), .A2(n684), .ZN(G66) );
  XOR2_X1 U736 ( .A(n686), .B(KEYINPUT121), .Z(n687) );
  NOR2_X1 U737 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U738 ( .A(KEYINPUT122), .B(n689), .Z(n696) );
  NAND2_X1 U739 ( .A1(G224), .A2(G953), .ZN(n690) );
  XNOR2_X1 U740 ( .A(n690), .B(KEYINPUT61), .ZN(n691) );
  XNOR2_X1 U741 ( .A(KEYINPUT120), .B(n691), .ZN(n692) );
  NAND2_X1 U742 ( .A1(G898), .A2(n692), .ZN(n694) );
  NAND2_X1 U743 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U744 ( .A(n696), .B(n695), .Z(G69) );
  XOR2_X1 U745 ( .A(n698), .B(n697), .Z(n704) );
  XOR2_X1 U746 ( .A(G227), .B(n704), .Z(n699) );
  XNOR2_X1 U747 ( .A(n699), .B(KEYINPUT123), .ZN(n700) );
  NAND2_X1 U748 ( .A1(n700), .A2(G900), .ZN(n701) );
  NAND2_X1 U749 ( .A1(G953), .A2(n701), .ZN(n702) );
  XNOR2_X1 U750 ( .A(n702), .B(KEYINPUT124), .ZN(n708) );
  XOR2_X1 U751 ( .A(n704), .B(n703), .Z(n706) );
  NAND2_X1 U752 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U753 ( .A1(n708), .A2(n707), .ZN(G72) );
  XNOR2_X1 U754 ( .A(n709), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U755 ( .A(G122), .B(KEYINPUT125), .Z(n710) );
  XNOR2_X1 U756 ( .A(n711), .B(n710), .ZN(G24) );
  XNOR2_X1 U757 ( .A(G110), .B(n712), .ZN(G12) );
  XNOR2_X1 U758 ( .A(G140), .B(KEYINPUT115), .ZN(n714) );
  XNOR2_X1 U759 ( .A(n714), .B(n713), .ZN(G42) );
  XNOR2_X1 U760 ( .A(n715), .B(G131), .ZN(G33) );
  XNOR2_X1 U761 ( .A(G134), .B(n716), .ZN(G36) );
  XOR2_X1 U762 ( .A(G137), .B(n717), .Z(n718) );
  XNOR2_X1 U763 ( .A(KEYINPUT127), .B(n718), .ZN(G39) );
endmodule

