//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT8), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(new_n214), .A3(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n254), .A2(new_n255), .A3(new_n213), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n254), .B2(new_n213), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n253), .A2(new_n258), .B1(new_n202), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  XOR2_X1   g0066(.A(new_n266), .B(KEYINPUT71), .Z(new_n267));
  NAND2_X1  g0067(.A1(new_n254), .A2(new_n213), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n254), .A2(new_n255), .A3(new_n213), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n267), .A2(new_n261), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n213), .ZN(new_n277));
  AND2_X1   g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(KEYINPUT67), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n291), .A2(new_n292), .A3(new_n283), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G77), .B2(new_n291), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n281), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n278), .A2(new_n279), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(new_n224), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT68), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n295), .A2(KEYINPUT68), .A3(new_n301), .ZN(new_n304));
  OAI21_X1  g0104(.A(G179), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n304), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G169), .A3(new_n302), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n274), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(G190), .B1(new_n303), .B2(new_n304), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(G200), .A3(new_n302), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n273), .B(KEYINPUT9), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n309), .A2(new_n310), .A3(new_n311), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n308), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n298), .B1(new_n300), .B2(new_n226), .ZN(new_n317));
  INV_X1    g0117(.A(new_n281), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G238), .A2(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n234), .B2(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n282), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G107), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n282), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G190), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT72), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G20), .A2(G77), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(new_n251), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n214), .A2(G33), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT15), .B(G87), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n331), .B1(new_n332), .B2(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n258), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n271), .A2(G77), .A3(new_n261), .A4(new_n265), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n262), .A2(new_n225), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n337), .A2(KEYINPUT73), .A3(new_n338), .A4(new_n339), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n324), .A2(G179), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n324), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT74), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n271), .A2(G68), .A3(new_n261), .A4(new_n265), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n260), .A2(G20), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n353), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n354), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n225), .B2(new_n334), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n258), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT11), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G232), .A2(G1698), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n224), .B2(G1698), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n282), .A2(new_n370), .B1(G33), .B2(G97), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n281), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n298), .B1(new_n300), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT75), .B(KEYINPUT13), .C1(new_n372), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n296), .A2(new_n297), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n299), .A2(new_n296), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(G238), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n378), .B(new_n379), .C1(new_n281), .C2(new_n371), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(new_n380), .A3(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n378), .B(KEYINPUT13), .C1(new_n281), .C2(new_n371), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT13), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n372), .B2(new_n374), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT77), .B1(new_n368), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n366), .B1(new_n358), .B2(new_n360), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n381), .A4(new_n385), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n382), .A2(new_n384), .A3(G169), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n392), .A2(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n375), .A2(new_n380), .A3(G179), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n392), .B2(KEYINPUT14), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n368), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n316), .A2(new_n352), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n271), .A2(new_n261), .A3(new_n265), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n249), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n262), .B2(new_n249), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT80), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n399), .B(new_n402), .C1(new_n262), .C2(new_n249), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G58), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n354), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n406), .A2(new_n201), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n287), .B2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n289), .A2(KEYINPUT78), .A3(G33), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n288), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n413), .B2(new_n214), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(KEYINPUT79), .A3(KEYINPUT7), .A4(new_n214), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n409), .B1(new_n419), .B2(G68), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n271), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n282), .B2(G20), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n427), .B2(new_n408), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n404), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n299), .A2(G232), .A3(new_n296), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT81), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n298), .B1(new_n431), .B2(KEYINPUT81), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT82), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT81), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n377), .A2(new_n436), .A3(G232), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT82), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n432), .A4(new_n298), .ZN(new_n439));
  MUX2_X1   g0239(.A(new_n292), .B(new_n224), .S(G1698), .Z(new_n440));
  OAI22_X1  g0240(.A1(new_n413), .A2(new_n440), .B1(new_n287), .B2(new_n218), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n318), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n435), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n348), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G179), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n430), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n419), .A2(G68), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n258), .A3(new_n429), .ZN(new_n449));
  INV_X1    g0249(.A(new_n404), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n328), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G190), .B2(new_n443), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n445), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n271), .B(new_n428), .C1(new_n420), .C2(KEYINPUT16), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n404), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n449), .A2(new_n450), .A3(new_n452), .A4(KEYINPUT17), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n446), .A2(new_n455), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n397), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT21), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n264), .A2(G33), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n261), .B(new_n464), .C1(new_n256), .C2(new_n257), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  INV_X1    g0266(.A(new_n260), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT86), .A2(G116), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT86), .A2(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT20), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n214), .C1(G33), .C2(new_n220), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n268), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n468), .A2(new_n469), .A3(new_n214), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT89), .B(new_n473), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n471), .A2(KEYINPUT20), .A3(new_n475), .A4(new_n268), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT86), .B(G116), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n268), .B(new_n475), .C1(new_n481), .C2(new_n214), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT89), .B1(new_n482), .B2(new_n473), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n291), .A2(G303), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G264), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n221), .B2(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(new_n411), .A3(new_n288), .A4(new_n412), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n281), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n492), .B(G274), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n299), .ZN(new_n497));
  INV_X1    g0297(.A(G270), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n463), .B1(new_n485), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n495), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n496), .A2(new_n299), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G270), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n489), .A2(new_n486), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n318), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(G179), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n500), .B2(new_n463), .ZN(new_n508));
  INV_X1    g0308(.A(new_n472), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n478), .A2(new_n479), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n483), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n490), .A2(new_n499), .A3(G190), .ZN(new_n513));
  AOI21_X1  g0313(.A(G200), .B1(new_n504), .B2(new_n506), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n485), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n501), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n271), .A2(G107), .A3(new_n261), .A4(new_n464), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n264), .A2(new_n322), .A3(G13), .A4(G20), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT90), .B(KEYINPUT25), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT91), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT91), .B1(new_n525), .B2(new_n518), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n518), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT92), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n517), .B2(new_n528), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n214), .B(G33), .C1(new_n468), .C2(new_n469), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n214), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n322), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n218), .A2(G20), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT22), .B1(new_n282), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT78), .B1(new_n289), .B2(G33), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n289), .A2(G33), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT22), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n218), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n214), .A3(new_n412), .A4(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n539), .A2(new_n542), .A3(new_n548), .A4(KEYINPUT24), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n258), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n538), .A2(new_n541), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT24), .B1(new_n551), .B2(new_n548), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n531), .A2(new_n532), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G257), .A2(G1698), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n219), .B2(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(new_n411), .A3(new_n288), .A4(new_n412), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G294), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n318), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n496), .A2(G264), .A3(new_n299), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n561), .A3(new_n495), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n328), .ZN(new_n563));
  INV_X1    g0363(.A(G190), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n281), .B1(new_n557), .B2(new_n556), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n502), .A3(new_n560), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n563), .A2(KEYINPUT93), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT93), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n568), .A3(new_n328), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n553), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n552), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n411), .A2(new_n412), .A3(new_n214), .A4(new_n288), .ZN(new_n572));
  INV_X1    g0372(.A(new_n547), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n574), .A2(new_n541), .A3(new_n538), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n271), .B1(new_n575), .B2(KEYINPUT24), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n517), .A2(new_n528), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT92), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n571), .A2(new_n576), .B1(new_n578), .B2(new_n530), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n560), .B1(new_n318), .B2(new_n558), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n348), .B1(new_n580), .B2(new_n495), .ZN(new_n581));
  INV_X1    g0381(.A(G179), .ZN(new_n582));
  NOR4_X1   g0382(.A1(new_n565), .A2(new_n560), .A3(new_n582), .A4(new_n502), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n516), .A2(new_n570), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n495), .B1(new_n497), .B2(new_n221), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n283), .A2(G244), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n413), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G250), .A2(G1698), .ZN(new_n592));
  NAND2_X1  g0392(.A1(KEYINPUT4), .A2(G244), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(G1698), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n282), .A2(new_n594), .B1(G33), .B2(G283), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(KEYINPUT84), .B(new_n588), .C1(new_n596), .C2(new_n281), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n281), .B1(new_n591), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n587), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n348), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n599), .A2(new_n587), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n582), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT6), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n605), .A2(new_n220), .A3(G107), .ZN(new_n606));
  XNOR2_X1  g0406(.A(G97), .B(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n608), .A2(new_n214), .B1(new_n225), .B2(new_n333), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n322), .B1(new_n423), .B2(new_n425), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n258), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n465), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G97), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n261), .A2(G97), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n602), .A2(new_n604), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n597), .A2(G190), .A3(new_n600), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n611), .A2(KEYINPUT83), .A3(new_n613), .A4(new_n615), .ZN(new_n621));
  INV_X1    g0421(.A(new_n603), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n465), .A2(new_n218), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(G33), .A2(G97), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT19), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n214), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(G87), .A2(G97), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n322), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(KEYINPUT87), .B(new_n628), .C1(new_n627), .C2(G20), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT87), .B1(new_n635), .B2(new_n628), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n572), .A2(new_n354), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n258), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n335), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n261), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n626), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n481), .A2(G33), .ZN(new_n644));
  NAND2_X1  g0444(.A1(G244), .A2(G1698), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n373), .B2(G1698), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n411), .A3(new_n288), .A4(new_n412), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n281), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  OAI221_X1 g0448(.A(G250), .B1(G1), .B2(new_n491), .C1(new_n276), .C2(new_n213), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n492), .A2(KEYINPUT85), .A3(G274), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n264), .A2(G45), .A3(G274), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT85), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(G200), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT88), .B1(new_n643), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n647), .A2(new_n644), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n318), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(G190), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n545), .A2(new_n214), .A3(G68), .A4(new_n412), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n628), .B1(new_n627), .B2(G20), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n633), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(new_n632), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n641), .B1(new_n667), .B2(new_n258), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n655), .A4(new_n626), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n657), .A2(new_n661), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n271), .A2(new_n261), .A3(new_n640), .A4(new_n464), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n639), .A2(new_n642), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n659), .A2(new_n660), .A3(new_n582), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n348), .B1(new_n648), .B2(new_n654), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n617), .A2(new_n624), .A3(new_n671), .A4(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n462), .A2(new_n586), .A3(new_n677), .ZN(G372));
  NAND4_X1  g0478(.A1(new_n668), .A2(new_n655), .A3(new_n626), .A4(new_n661), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT93), .B1(new_n566), .B2(G200), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n566), .A2(new_n564), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n569), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n680), .B1(new_n579), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n501), .B(new_n512), .C1(new_n579), .C2(new_n584), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n617), .A3(new_n685), .A4(new_n624), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n670), .A2(new_n661), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n665), .A2(new_n633), .B1(new_n629), .B2(new_n631), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n271), .B1(new_n688), .B2(new_n662), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n689), .A2(new_n625), .A3(new_n641), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n669), .B1(new_n690), .B2(new_n655), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n676), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT26), .B1(new_n692), .B2(new_n617), .ZN(new_n693));
  INV_X1    g0493(.A(new_n680), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n601), .A2(new_n348), .B1(new_n582), .B2(new_n603), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n619), .A2(new_n621), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n676), .B(KEYINPUT94), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n686), .A2(new_n693), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n462), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n446), .A2(new_n459), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n350), .B1(new_n387), .B2(new_n390), .ZN(new_n703));
  INV_X1    g0503(.A(new_n396), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n455), .B(new_n460), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n313), .A2(new_n315), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n308), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(new_n708), .ZN(G369));
  INV_X1    g0509(.A(new_n585), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n467), .A2(KEYINPUT27), .A3(G20), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT27), .B1(new_n467), .B2(G20), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G343), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n683), .A2(new_n579), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n579), .B2(new_n715), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n710), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n501), .A2(new_n512), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n716), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT95), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(KEYINPUT95), .A3(new_n718), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n721), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n717), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n485), .A2(new_n715), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n722), .B2(new_n515), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n722), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n728), .A2(new_n737), .ZN(G399));
  INV_X1    g0538(.A(new_n208), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G41), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G1), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n630), .A2(new_n322), .A3(new_n466), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n743), .B1(new_n211), .B2(new_n741), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  INV_X1    g0545(.A(G330), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n648), .A2(new_n654), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n747), .A2(new_n580), .ZN(new_n748));
  INV_X1    g0548(.A(new_n507), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n600), .A4(new_n597), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(G179), .B1(new_n504), .B2(new_n506), .ZN(new_n753));
  INV_X1    g0553(.A(new_n747), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n622), .A2(new_n753), .A3(new_n562), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n750), .B2(new_n751), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n716), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n677), .A2(new_n586), .A3(new_n715), .ZN(new_n761));
  OAI211_X1 g0561(.A(KEYINPUT31), .B(new_n716), .C1(new_n752), .C2(new_n756), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n746), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n700), .A2(new_n715), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT29), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n617), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n697), .A3(new_n676), .A4(new_n671), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT26), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n769), .A2(new_n686), .A3(new_n699), .A4(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(KEYINPUT29), .A3(new_n715), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n764), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n745), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n259), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n742), .B1(G45), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n735), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n734), .A2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n734), .A2(G20), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n739), .A2(new_n291), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G355), .B1(new_n466), .B2(new_n739), .ZN(new_n787));
  INV_X1    g0587(.A(new_n413), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n739), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n212), .A2(G45), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n242), .B2(G45), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n783), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n213), .B1(G20), .B2(new_n348), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n214), .A2(new_n564), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n582), .A2(G200), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n291), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n214), .A2(G190), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n328), .A2(G179), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G179), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G283), .A2(new_n807), .B1(new_n810), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n798), .A2(new_n805), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n582), .A2(new_n328), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(new_n798), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n811), .B1(new_n812), .B2(new_n813), .C1(new_n814), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n808), .A2(G190), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G20), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n803), .B(new_n818), .C1(G294), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT100), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n815), .A2(new_n822), .A3(new_n804), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n815), .B2(new_n804), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n804), .A2(new_n799), .A3(KEYINPUT98), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT98), .B1(new_n804), .B2(new_n799), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n826), .A2(new_n827), .B1(new_n831), .B2(G311), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n813), .A2(new_n218), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n291), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  INV_X1    g0635(.A(new_n820), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n220), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G107), .A2(new_n807), .B1(new_n816), .B2(G50), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n405), .B2(new_n801), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n810), .A2(G159), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT32), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n825), .A2(new_n354), .B1(new_n830), .B2(new_n225), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n821), .A2(new_n832), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n795), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n797), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n777), .B1(new_n784), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n781), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NAND2_X1  g0651(.A1(new_n846), .A2(new_n783), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(G77), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n778), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n826), .A2(G283), .B1(G303), .B2(new_n816), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n470), .B2(new_n830), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT102), .Z(new_n857));
  OAI21_X1  g0657(.A(new_n291), .B1(new_n813), .B2(new_n322), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n807), .A2(G87), .ZN(new_n860));
  INV_X1    g0660(.A(G311), .ZN(new_n861));
  INV_X1    g0661(.A(G294), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n809), .C1(new_n801), .C2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n859), .A2(new_n863), .A3(new_n837), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n816), .B1(new_n800), .B2(G143), .ZN(new_n865));
  INV_X1    g0665(.A(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G150), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n865), .B1(new_n830), .B2(new_n866), .C1(new_n825), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT34), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n806), .A2(new_n354), .ZN(new_n870));
  INV_X1    g0670(.A(new_n813), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(G50), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n809), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n413), .B(new_n874), .C1(G58), .C2(new_n820), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n857), .A2(new_n864), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n350), .A2(new_n716), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n715), .B1(new_n342), .B2(new_n343), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n330), .B2(new_n345), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n880), .B2(new_n350), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n854), .B1(new_n846), .B2(new_n876), .C1(new_n881), .C2(new_n783), .ZN(new_n882));
  INV_X1    g0682(.A(new_n877), .ZN(new_n883));
  INV_X1    g0683(.A(new_n350), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n765), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n700), .A2(new_n715), .A3(new_n881), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n764), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n778), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n764), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT104), .Z(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(G384));
  INV_X1    g0693(.A(new_n608), .ZN(new_n894));
  OAI211_X1 g0694(.A(G116), .B(new_n215), .C1(new_n894), .C2(KEYINPUT35), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(KEYINPUT35), .B2(new_n894), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n406), .A2(new_n211), .A3(new_n225), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT105), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n898), .A2(new_n899), .B1(new_n202), .B2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n264), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n761), .A2(new_n762), .A3(new_n759), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n391), .A2(new_n396), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n388), .A2(new_n715), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n391), .B(new_n396), .C1(new_n388), .C2(new_n715), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n885), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n904), .A2(new_n909), .A3(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT16), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n354), .B1(new_n417), .B2(new_n418), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n912), .B2(new_n409), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n404), .B1(new_n421), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n453), .B1(new_n914), .B2(new_n713), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n445), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n449), .A2(new_n450), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n456), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n714), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n453), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n914), .A2(new_n713), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n461), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n453), .B1(new_n430), .B2(new_n445), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n430), .A2(new_n713), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT37), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n461), .A2(new_n928), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n910), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n910), .B(KEYINPUT107), .C1(new_n926), .C2(new_n932), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n904), .A2(new_n909), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n923), .B2(new_n925), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n462), .A2(new_n904), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n941), .B(new_n942), .Z(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n746), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n396), .A2(new_n716), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT39), .B1(new_n926), .B2(new_n939), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n922), .A2(new_n929), .B1(new_n461), .B2(new_n928), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n949), .C1(KEYINPUT38), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n907), .A2(new_n908), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n887), .B2(new_n883), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n926), .B2(new_n939), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n702), .A2(new_n714), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n462), .A2(new_n767), .A3(new_n773), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n462), .A2(new_n773), .A3(KEYINPUT106), .A4(new_n767), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n708), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n959), .B(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n944), .A2(new_n965), .B1(new_n264), .B2(new_n776), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n944), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n903), .B1(new_n966), .B2(new_n967), .ZN(G367));
  NOR2_X1   g0768(.A1(new_n690), .A2(new_n715), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n699), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n694), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n794), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT46), .B1(new_n871), .B2(new_n481), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n413), .B1(new_n801), .B2(new_n812), .C1(new_n861), .C2(new_n817), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G107), .C2(new_n820), .ZN(new_n975));
  INV_X1    g0775(.A(G283), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n830), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n871), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n810), .A2(G317), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n220), .C2(new_n806), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(G294), .C2(new_n826), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n282), .B1(new_n806), .B2(new_n225), .C1(new_n836), .C2(new_n354), .ZN(new_n982));
  INV_X1    g0782(.A(G143), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n817), .A2(new_n983), .B1(new_n801), .B2(new_n867), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n813), .A2(new_n405), .B1(new_n809), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n826), .A2(G159), .B1(new_n831), .B2(G50), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n975), .A2(new_n981), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n846), .B1(new_n989), .B2(KEYINPUT47), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT47), .B2(new_n989), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n796), .B1(new_n208), .B2(new_n335), .C1(new_n790), .C2(new_n238), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n972), .A2(new_n777), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n724), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n715), .B1(new_n619), .B2(new_n621), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n617), .A3(new_n624), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n695), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT42), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n768), .B1(new_n999), .B2(new_n585), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n716), .B1(new_n1002), .B2(KEYINPUT108), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(KEYINPUT108), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(KEYINPUT42), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1004), .A2(KEYINPUT109), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT109), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT110), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n1001), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT43), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n971), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n971), .A2(new_n1012), .ZN(new_n1014));
  AND4_X1   g0814(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n999), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n737), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n776), .A2(G45), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(G1), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n726), .A2(new_n727), .A3(new_n1017), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n726), .A2(new_n727), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1029), .A2(KEYINPUT111), .A3(KEYINPUT44), .A4(new_n1017), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT112), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1025), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT111), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n728), .A2(new_n999), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT45), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n736), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n737), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n730), .A2(new_n723), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n994), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(new_n735), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n774), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n774), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n740), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1024), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n993), .B1(new_n1022), .B2(new_n1049), .ZN(G387));
  AOI22_X1  g0850(.A1(G322), .A2(new_n816), .B1(new_n800), .B2(G317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n830), .B2(new_n812), .C1(new_n825), .C2(new_n861), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n871), .A2(G294), .B1(new_n820), .B2(G283), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT49), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n413), .B1(new_n809), .B2(new_n814), .C1(new_n470), .C2(new_n806), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n871), .A2(G77), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n867), .B2(new_n809), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G159), .B2(new_n816), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n831), .A2(G68), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n826), .A2(new_n249), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n836), .A2(new_n335), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n801), .A2(new_n202), .B1(new_n806), .B2(new_n220), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1068), .A2(new_n413), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n795), .B1(new_n1062), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n790), .B1(new_n235), .B2(G45), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n743), .B2(new_n786), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n332), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n202), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n491), .B1(new_n354), .B2(new_n225), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n743), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1074), .A2(new_n1079), .B1(G107), .B2(new_n208), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n796), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1072), .A2(new_n1081), .A3(new_n777), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n731), .B2(new_n794), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1044), .B2(new_n1024), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1044), .A2(new_n774), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1044), .A2(new_n774), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n740), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(G393));
  NAND3_X1  g0889(.A1(new_n1040), .A2(new_n1041), .A3(new_n1024), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1017), .A2(new_n794), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n860), .B1(new_n354), .B2(new_n813), .C1(new_n983), .C2(new_n809), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n413), .B(new_n1092), .C1(G77), .C2(new_n820), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n826), .A2(G50), .B1(new_n831), .B2(new_n1075), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G150), .A2(new_n816), .B1(new_n800), .B2(G159), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G283), .A2(new_n871), .B1(new_n810), .B2(G322), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n291), .C1(new_n322), .C2(new_n806), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT115), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G317), .A2(new_n816), .B1(new_n800), .B2(G311), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n862), .C2(new_n830), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n825), .A2(new_n812), .B1(new_n470), .B2(new_n836), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT116), .Z(new_n1106));
  OAI21_X1  g0906(.A(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n795), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n796), .B1(new_n220), .B2(new_n208), .C1(new_n790), .C2(new_n245), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1091), .A2(new_n777), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1090), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1045), .A2(new_n740), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1087), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G390));
  NAND2_X1  g0916(.A1(new_n887), .A2(new_n883), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n953), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n946), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n947), .A2(new_n1119), .A3(new_n951), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n948), .B1(new_n950), .B2(KEYINPUT38), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n880), .A2(new_n350), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n772), .A2(new_n715), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n883), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n953), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n945), .B(KEYINPUT117), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n764), .A2(new_n909), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1120), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n904), .A2(new_n953), .A3(G330), .A4(new_n881), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT118), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1131), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n953), .B1(new_n764), .B2(new_n881), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1117), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n904), .A2(G330), .A3(new_n881), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n954), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1128), .A2(new_n883), .A3(new_n1123), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n462), .A2(G330), .A3(new_n904), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n962), .A2(new_n708), .A3(new_n963), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n741), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1133), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n947), .A2(new_n782), .A3(new_n951), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n777), .B1(new_n249), .B2(new_n852), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n826), .A2(G107), .B1(new_n831), .B2(G97), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n870), .B1(G294), .B2(new_n810), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G283), .A2(new_n816), .B1(new_n800), .B2(G116), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n282), .B(new_n833), .C1(G77), .C2(new_n820), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n813), .A2(new_n867), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n985), .B2(new_n825), .C1(new_n830), .C2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G50), .A2(new_n807), .B1(new_n816), .B2(G128), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n800), .A2(G132), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n820), .A2(G159), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n291), .B1(new_n810), .B2(G125), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1155), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1150), .B1(new_n1165), .B2(new_n795), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1149), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1024), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1134), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1148), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n951), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n923), .A2(new_n925), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT38), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n949), .B1(new_n1176), .B2(new_n948), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n945), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n958), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1180), .A2(new_n941), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n940), .A2(new_n937), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n936), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT107), .B1(new_n1121), .B2(new_n910), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G330), .B(new_n1182), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n959), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1189));
  NAND2_X1  g0989(.A1(new_n316), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n316), .A2(new_n1189), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n273), .A2(new_n714), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT55), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1193), .B(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1188), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT121), .B1(new_n941), .B2(G330), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1181), .B(new_n1187), .C1(new_n1200), .C2(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1143), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1172), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(KEYINPUT57), .B(new_n1203), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n740), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(new_n1024), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1197), .A2(new_n782), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n777), .B1(G50), .B2(new_n852), .ZN(new_n1211));
  INV_X1    g1011(.A(G41), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G50), .B1(new_n287), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n788), .B2(G41), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT119), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1063), .B1(new_n817), .B2(new_n466), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n807), .A2(G58), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n976), .B2(new_n809), .C1(new_n801), .C2(new_n322), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G68), .C2(new_n820), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G41), .B(new_n788), .C1(new_n831), .C2(new_n640), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n220), .C2(new_n825), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1215), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n816), .A2(G125), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1224), .B1(new_n813), .B2(new_n1158), .C1(new_n801), .C2(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n825), .A2(new_n873), .B1(new_n830), .B2(new_n985), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(G150), .C2(new_n820), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n287), .B(new_n1212), .C1(new_n806), .C2(new_n866), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G124), .B2(new_n810), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT59), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1230), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1211), .B1(new_n1235), .B2(new_n795), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1210), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1209), .A2(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1208), .A2(KEYINPUT122), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1238), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1207), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1239), .A2(new_n1242), .ZN(G375));
  OAI221_X1 g1043(.A(new_n1217), .B1(new_n1225), .B2(new_n809), .C1(new_n866), .C2(new_n813), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n413), .B(new_n1244), .C1(G50), .C2(new_n820), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n817), .A2(new_n873), .B1(new_n801), .B2(new_n985), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1158), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n826), .B2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n831), .A2(G150), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1245), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n282), .B(new_n1069), .C1(G77), .C2(new_n807), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n816), .A2(G294), .B1(new_n810), .B2(G303), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n826), .A2(new_n481), .B1(new_n831), .B2(G107), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G97), .A2(new_n871), .B1(new_n800), .B2(G283), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n777), .B1(G68), .B2(new_n852), .C1(new_n1258), .C2(new_n846), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n954), .B2(new_n782), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1141), .B2(new_n1024), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1168), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT125), .B1(new_n1264), .B2(new_n1260), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1137), .A2(new_n1143), .A3(new_n1140), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1047), .B(KEYINPUT123), .Z(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1145), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G381));
  OAI21_X1  g1071(.A(new_n1170), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1047), .B1(new_n1045), .B2(new_n774), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1020), .B(new_n1021), .C1(new_n1274), .C2(new_n1024), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1275), .A2(new_n993), .A3(new_n1115), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1276), .A3(new_n1277), .ZN(G407));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G343), .C2(new_n1272), .ZN(G409));
  XNOR2_X1  g1079(.A(G393), .B(new_n850), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1115), .B1(new_n1275), .B2(new_n993), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1276), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G387), .A2(G390), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1275), .A2(new_n993), .A3(new_n1115), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1280), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1207), .A2(G378), .A3(new_n1241), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1268), .B(new_n1203), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1170), .B1(new_n1238), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(G343), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G213), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n741), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1297));
  OAI211_X1 g1097(.A(KEYINPUT126), .B(new_n1295), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1266), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1267), .B(KEYINPUT60), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1300), .B2(new_n1295), .ZN(new_n1301));
  OAI21_X1  g1101(.A(G384), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1305), .A2(new_n892), .A3(new_n1266), .A4(new_n1298), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1291), .A2(new_n1292), .A3(new_n1294), .A4(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1288), .A2(new_n1290), .B1(G213), .B2(new_n1293), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1293), .A2(G213), .A3(G2897), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1302), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1308), .B(new_n1309), .C1(new_n1310), .C2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1292), .B1(new_n1310), .B2(new_n1307), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1287), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT63), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1307), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1287), .A2(KEYINPUT61), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1317), .A2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(new_n1287), .A2(new_n1307), .ZN(new_n1325));
  OAI21_X1  g1125(.A(G378), .B1(new_n1208), .B2(new_n1238), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1282), .A2(new_n1286), .A3(new_n1306), .A4(new_n1302), .ZN(new_n1327));
  AND4_X1   g1127(.A1(new_n1272), .A2(new_n1325), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n1325), .A2(new_n1327), .B1(new_n1272), .B2(new_n1326), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


