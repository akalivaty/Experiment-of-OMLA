//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n228), .A2(new_n213), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n216), .B(new_n222), .C1(new_n223), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n223), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G107), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT25), .B1(new_n253), .B2(new_n254), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n210), .A2(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n252), .A2(new_n258), .A3(new_n220), .A4(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT24), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n254), .A2(KEYINPUT23), .A3(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT23), .B1(new_n254), .B2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G116), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n263), .A2(new_n264), .B1(G20), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT22), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n211), .A3(G87), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n262), .B1(new_n270), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n270), .A2(new_n262), .A3(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n259), .A2(new_n220), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n261), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT84), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n271), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n268), .B2(new_n275), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G257), .A2(G1698), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G250), .ZN(new_n292));
  XOR2_X1   g0092(.A(KEYINPUT85), .B(G294), .Z(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n278), .A2(KEYINPUT84), .A3(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n290), .A2(new_n292), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT86), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  INV_X1    g0101(.A(new_n220), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT76), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n210), .B(G45), .C1(new_n305), .C2(KEYINPUT5), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT75), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G1), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT5), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G41), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n308), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n311), .A3(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n307), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n306), .A3(new_n319), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n322), .A2(G264), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n300), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n327));
  OAI21_X1  g0127(.A(G169), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n297), .A2(new_n299), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(new_n325), .A3(G179), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n285), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n282), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n284), .B1(new_n332), .B2(new_n280), .ZN(new_n333));
  INV_X1    g0133(.A(new_n261), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(KEYINPUT86), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n300), .A4(new_n325), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(new_n325), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n322), .A2(G257), .A3(new_n323), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT77), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT77), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n322), .A2(new_n346), .A3(G257), .A4(new_n323), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n307), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT76), .B1(new_n318), .B2(new_n319), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n278), .A2(G244), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT4), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n356), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G283), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G244), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n276), .B2(new_n277), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT4), .B1(new_n368), .B2(new_n356), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT74), .B1(new_n369), .B2(new_n363), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n299), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n352), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n355), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n354), .B(new_n321), .C1(new_n345), .C2(new_n347), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT78), .B1(new_n348), .B2(new_n352), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(G190), .A3(new_n372), .ZN(new_n379));
  INV_X1    g0179(.A(new_n284), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G20), .A2(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G77), .ZN(new_n382));
  XOR2_X1   g0182(.A(new_n382), .B(KEYINPUT72), .Z(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(G97), .A3(new_n254), .ZN(new_n385));
  XOR2_X1   g0185(.A(G97), .B(G107), .Z(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n383), .B1(new_n387), .B2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n272), .A2(new_n274), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n389), .B2(new_n211), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n391), .B(G20), .C1(new_n272), .C2(new_n274), .ZN(new_n392));
  OAI21_X1  g0192(.A(G107), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n380), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G97), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n253), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n260), .B2(new_n395), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n375), .A2(new_n379), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n323), .B1(new_n366), .B2(new_n370), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(G179), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n398), .B1(new_n378), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n374), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n278), .A2(G238), .A3(new_n356), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(new_n265), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n299), .ZN(new_n409));
  INV_X1    g0209(.A(G250), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n312), .B2(G1), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n210), .A2(new_n301), .A3(G45), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n323), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n323), .A2(new_n411), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n340), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n337), .B(new_n417), .C1(new_n408), .C2(new_n299), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI211_X1 g0221(.A(G20), .B(new_n246), .C1(new_n276), .C2(new_n277), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n211), .A2(G33), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n423), .A2(KEYINPUT19), .A3(new_n395), .ZN(new_n424));
  INV_X1    g0224(.A(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n207), .A2(new_n425), .B1(new_n426), .B2(new_n211), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(KEYINPUT19), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT80), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n278), .A2(new_n211), .A3(G68), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT19), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n431), .B(new_n432), .C1(new_n434), .C2(new_n424), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n435), .A3(new_n284), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n253), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n260), .A2(new_n425), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n265), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n291), .B2(G238), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n323), .B1(new_n442), .B2(new_n406), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n443), .B2(new_n417), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n409), .A2(G179), .A3(new_n418), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n260), .A2(new_n437), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n436), .A2(new_n438), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n421), .A2(new_n440), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n343), .A2(new_n399), .A3(new_n405), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n268), .A2(G222), .A3(new_n356), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n389), .A2(new_n356), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(G223), .B1(G77), .B2(new_n389), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n323), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G1), .B1(new_n305), .B2(new_n312), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n323), .A3(G274), .ZN(new_n458));
  INV_X1    g0258(.A(G226), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n323), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G190), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n204), .A2(new_n211), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT67), .A2(G58), .ZN(new_n466));
  XOR2_X1   g0266(.A(new_n466), .B(KEYINPUT8), .Z(new_n467));
  INV_X1    g0267(.A(G150), .ZN(new_n468));
  INV_X1    g0268(.A(new_n381), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n467), .A2(new_n423), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n284), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n252), .A2(G50), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n284), .B1(new_n210), .B2(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(G50), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT9), .ZN(new_n476));
  OAI21_X1  g0276(.A(G200), .B1(new_n456), .B2(new_n462), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n474), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT9), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n464), .A2(new_n476), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT10), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n478), .B(KEYINPUT9), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT10), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n477), .A4(new_n464), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G179), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n463), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n403), .B1(new_n456), .B2(new_n462), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n478), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n381), .A2(G50), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT69), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n423), .A2(new_n205), .B1(new_n211), .B2(G68), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n284), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT11), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n500));
  AOI22_X1  g0300(.A1(G68), .A2(new_n473), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT14), .ZN(new_n503));
  INV_X1    g0303(.A(new_n458), .ZN(new_n504));
  INV_X1    g0304(.A(new_n461), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(G238), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT13), .ZN(new_n507));
  INV_X1    g0307(.A(G232), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G1698), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G226), .B2(G1698), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n426), .B1(new_n510), .B2(new_n389), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n299), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n506), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n507), .B1(new_n506), .B2(new_n512), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n503), .B(G169), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n487), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n503), .B1(new_n516), .B2(G169), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n502), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(G200), .ZN(new_n520));
  INV_X1    g0320(.A(new_n502), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n337), .C2(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n491), .B1(new_n524), .B2(KEYINPUT70), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G87), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G223), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n459), .B2(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n288), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n299), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n505), .A2(G232), .B1(new_n304), .B2(new_n457), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n403), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n458), .B1(new_n508), .B2(new_n461), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n487), .B(new_n534), .C1(new_n530), .C2(new_n299), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G58), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n246), .ZN(new_n538));
  OAI21_X1  g0338(.A(G20), .B1(new_n538), .B2(new_n201), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n381), .A2(G159), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n391), .B1(new_n288), .B2(new_n211), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n276), .A2(new_n391), .A3(new_n211), .A4(new_n277), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G68), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT16), .B(new_n542), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n391), .B1(new_n268), .B2(G20), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n246), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(new_n541), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n284), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n467), .A2(new_n473), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n252), .B2(new_n467), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n536), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT18), .ZN(new_n558));
  OAI21_X1  g0358(.A(G68), .B1(new_n390), .B2(new_n392), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n542), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n380), .B1(new_n560), .B2(new_n547), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n554), .B1(new_n561), .B2(new_n546), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n278), .A2(new_n528), .B1(G33), .B2(G87), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n337), .B(new_n532), .C1(new_n563), .C2(new_n323), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n534), .B1(new_n530), .B2(new_n299), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(KEYINPUT17), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT18), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n536), .A2(new_n556), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n552), .A2(new_n566), .A3(new_n555), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n558), .A2(new_n567), .A3(new_n569), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n473), .A2(G77), .ZN(new_n575));
  XNOR2_X1  g0375(.A(KEYINPUT8), .B(G58), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n469), .B1(new_n211), .B2(new_n205), .ZN(new_n577));
  INV_X1    g0377(.A(new_n437), .ZN(new_n578));
  INV_X1    g0378(.A(new_n423), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI221_X1 g0380(.A(new_n575), .B1(G77), .B2(new_n252), .C1(new_n580), .C2(new_n380), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n454), .A2(G238), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n268), .A2(G232), .A3(new_n356), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n254), .C2(new_n268), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n299), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n504), .B1(G244), .B2(new_n505), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n581), .B1(new_n587), .B2(G200), .ZN(new_n588));
  INV_X1    g0388(.A(new_n587), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n589), .A2(KEYINPUT68), .A3(G190), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT68), .B1(new_n589), .B2(G190), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n581), .B1(new_n589), .B2(G169), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n587), .A2(G179), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT70), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n523), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n525), .A2(new_n574), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n260), .A2(KEYINPUT82), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT82), .B1(new_n260), .B2(new_n600), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n253), .A2(new_n600), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n362), .B(new_n211), .C1(G33), .C2(new_n395), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(G20), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n284), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n605), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(new_n604), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(G257), .A2(G1698), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(G264), .B2(new_n356), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n277), .B2(new_n276), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n268), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n299), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n322), .A2(G270), .A3(new_n323), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n352), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(KEYINPUT21), .A3(G169), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n352), .A2(G179), .A3(new_n619), .A4(new_n620), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n613), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n612), .A3(G169), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT83), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n629), .A3(new_n626), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n612), .B1(new_n621), .B2(G200), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n337), .B2(new_n621), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n451), .A2(new_n599), .A3(new_n631), .A4(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n446), .A2(new_n449), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n402), .A2(new_n404), .A3(new_n450), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n402), .A2(new_n404), .A3(new_n450), .A4(KEYINPUT26), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n398), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n376), .A2(new_n377), .A3(new_n400), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(G190), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n375), .B1(new_n404), .B2(new_n402), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n328), .A2(new_n330), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n335), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n342), .B1(new_n647), .B2(new_n631), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n648), .A3(new_n450), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n599), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n558), .A2(new_n569), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n595), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n522), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n519), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n567), .A2(new_n572), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n486), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n490), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n651), .A2(new_n660), .ZN(G369));
  NAND2_X1  g0461(.A1(new_n622), .A2(new_n623), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n612), .ZN(new_n663));
  INV_X1    g0463(.A(new_n630), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n629), .B1(new_n625), .B2(new_n626), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(G343), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n343), .A2(new_n666), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n331), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT88), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(KEYINPUT88), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n663), .B(new_n633), .C1(new_n664), .C2(new_n665), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n613), .A2(new_n676), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n666), .A2(new_n686), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n343), .B1(new_n285), .B2(new_n676), .ZN(new_n690));
  INV_X1    g0490(.A(new_n676), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n331), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n683), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT89), .Z(G399));
  INV_X1    g0496(.A(new_n214), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n218), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n650), .B2(new_n676), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI211_X1 g0506(.A(KEYINPUT29), .B(new_n691), .C1(new_n641), .C2(new_n649), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n623), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n443), .A2(new_n417), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n324), .B1(new_n297), .B2(new_n299), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n643), .A2(KEYINPUT30), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n374), .B2(new_n713), .ZN(new_n717));
  INV_X1    g0517(.A(new_n711), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n621), .A2(new_n487), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n374), .A2(new_n339), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n691), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n685), .A2(new_n691), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n645), .A2(new_n725), .A3(new_n343), .A4(new_n450), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n676), .A2(new_n723), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n717), .A2(new_n720), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  INV_X1    g0531(.A(new_n715), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n730), .B2(KEYINPUT90), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(G330), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n709), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n703), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(KEYINPUT91), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n689), .B(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n211), .A2(G13), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n210), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n698), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n687), .A2(new_n688), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n740), .B(new_n745), .C1(G330), .C2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n744), .B(KEYINPUT92), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n220), .B1(G20), .B2(new_n403), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n211), .A2(new_n487), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G200), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT95), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n337), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(G190), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G50), .A2(new_n756), .B1(new_n757), .B2(G68), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n211), .A2(G179), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n759), .A2(new_n337), .A3(G200), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(KEYINPUT32), .B1(new_n254), .B2(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n211), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(G97), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n752), .A2(new_n760), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n268), .B1(new_n771), .B2(new_n205), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n752), .A2(G190), .A3(new_n340), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G58), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n764), .A2(KEYINPUT32), .B1(new_n777), .B2(G87), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n758), .A2(new_n770), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT96), .B(G326), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n757), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  INV_X1    g0584(.A(G329), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n771), .A2(new_n784), .B1(new_n761), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n268), .B(new_n786), .C1(G322), .C2(new_n774), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n788), .A2(new_n765), .B1(new_n776), .B2(new_n617), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n293), .B2(new_n769), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n781), .A2(new_n783), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n751), .B1(new_n779), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n750), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n697), .A2(new_n389), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n600), .B2(new_n697), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n697), .A2(new_n278), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n312), .B2(new_n219), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n312), .B2(new_n250), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n749), .B(new_n792), .C1(new_n798), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n746), .B2(new_n796), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n747), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n750), .A2(new_n793), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n749), .B1(new_n205), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n595), .A2(new_n691), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n581), .A2(new_n691), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n592), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(new_n595), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n771), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n774), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(new_n757), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  INV_X1    g0620(.A(new_n756), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n818), .B1(new_n819), .B2(new_n468), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n768), .A2(new_n537), .B1(new_n776), .B2(new_n202), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n278), .B1(new_n827), .B2(new_n761), .ZN(new_n828));
  INV_X1    g0628(.A(new_n765), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(G68), .C2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n824), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n768), .A2(new_n395), .B1(new_n773), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT97), .Z(new_n834));
  OAI22_X1  g0634(.A1(new_n425), .A2(new_n765), .B1(new_n776), .B2(new_n254), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n389), .B1(new_n761), .B2(new_n784), .C1(new_n600), .C2(new_n771), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n757), .C2(G283), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n617), .B2(new_n821), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n831), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT98), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n750), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n812), .B1(new_n794), .B2(new_n816), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n650), .A2(new_n676), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n815), .A2(new_n595), .ZN(new_n847));
  INV_X1    g0647(.A(new_n813), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n592), .A2(new_n595), .A3(new_n676), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n641), .B2(new_n649), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n745), .B1(new_n855), .B2(new_n736), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(new_n735), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(G384));
  OR2_X1    g0658(.A1(new_n387), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n387), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(G116), .A3(new_n221), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n218), .A2(new_n205), .A3(new_n538), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n210), .B(G13), .C1(new_n864), .C2(new_n245), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n709), .A2(KEYINPUT105), .A3(new_n599), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT105), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n705), .A2(new_n707), .ZN(new_n869));
  INV_X1    g0669(.A(new_n599), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n660), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n653), .A2(new_n670), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n502), .A2(new_n691), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n519), .A2(new_n522), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n519), .B2(new_n522), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n852), .B2(new_n813), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n546), .A2(new_n284), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT7), .B1(new_n278), .B2(G20), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G68), .A3(new_n544), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT16), .B1(new_n882), .B2(new_n542), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n555), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n536), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n671), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n570), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT101), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT37), .B1(new_n556), .B2(new_n671), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(new_n557), .A3(new_n570), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n892), .A2(new_n893), .B1(new_n574), .B2(new_n886), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n891), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n886), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n573), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n894), .A2(new_n895), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n873), .B1(new_n879), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT102), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n873), .C1(new_n879), .C2(new_n902), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n562), .A2(new_n670), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n573), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n533), .A2(new_n535), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n570), .B1(new_n562), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n557), .A2(KEYINPUT103), .A3(new_n570), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n909), .B1(new_n562), .B2(new_n670), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n890), .A2(KEYINPUT104), .A3(new_n557), .A4(new_n570), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n908), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n895), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n901), .B1(new_n892), .B2(new_n893), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT39), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(KEYINPUT39), .B2(new_n902), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n519), .A2(new_n691), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n904), .A2(new_n906), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n872), .B(new_n929), .Z(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n728), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT106), .B1(new_n721), .B2(new_n728), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n724), .B(new_n726), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n877), .A2(new_n849), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n931), .B1(new_n936), .B2(new_n902), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n816), .B1(new_n875), .B2(new_n876), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n451), .A2(new_n725), .B1(new_n723), .B2(new_n722), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n721), .A2(new_n728), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n728), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n938), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n931), .B1(new_n922), .B2(new_n923), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n599), .A2(new_n934), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(G330), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n930), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT108), .Z(new_n954));
  OAI22_X1  g0754(.A1(new_n930), .A2(new_n952), .B1(new_n210), .B2(new_n741), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n866), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OR2_X1    g0759(.A1(new_n440), .A2(new_n676), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n450), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n960), .A2(new_n635), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n797), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n798), .B1(new_n214), .B2(new_n437), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n803), .A2(new_n240), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n748), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G143), .A2(new_n756), .B1(new_n757), .B2(G159), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n771), .A2(new_n202), .B1(new_n761), .B2(new_n820), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n389), .B(new_n972), .C1(G150), .C2(new_n774), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n765), .A2(new_n205), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n768), .A2(new_n246), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(G58), .C2(new_n777), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n776), .B2(new_n600), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT112), .ZN(new_n980));
  INV_X1    g0780(.A(new_n293), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n819), .B2(new_n981), .C1(new_n784), .C2(new_n821), .ZN(new_n982));
  INV_X1    g0782(.A(new_n761), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n774), .A2(G303), .B1(new_n983), .B2(G317), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n788), .B2(new_n771), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n288), .B1(new_n395), .B2(new_n765), .C1(new_n254), .C2(new_n768), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n776), .A2(new_n978), .A3(new_n600), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n970), .B1(new_n990), .B2(new_n750), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n967), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n737), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n642), .A2(new_n691), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n645), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n405), .B2(new_n676), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n683), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n405), .A2(new_n676), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n645), .B2(new_n995), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n681), .A2(new_n1000), .A3(KEYINPUT44), .A4(new_n682), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n677), .A2(KEYINPUT88), .A3(new_n678), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT88), .B1(new_n677), .B2(new_n678), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n683), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1002), .A2(new_n1009), .A3(new_n694), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n694), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n690), .B(new_n692), .C1(new_n631), .C2(new_n691), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1013), .A2(new_n689), .A3(new_n677), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n677), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n740), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1016), .A2(new_n735), .A3(new_n869), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n993), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n698), .B(KEYINPUT41), .Z(new_n1019));
  OAI21_X1  g0819(.A(new_n742), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n399), .A2(new_n331), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n405), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n676), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1000), .A2(new_n677), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT42), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT43), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n966), .B2(KEYINPUT110), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1028), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n694), .A2(new_n1000), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1032), .B(new_n1023), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT111), .B1(new_n1020), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n694), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1002), .A2(new_n1009), .A3(new_n694), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1017), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1019), .B1(new_n1047), .B2(new_n737), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1041), .B(KEYINPUT111), .C1(new_n1048), .C2(new_n743), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n992), .B1(new_n1042), .B2(new_n1050), .ZN(G387));
  AOI21_X1  g0851(.A(new_n278), .B1(new_n983), .B2(new_n780), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n981), .A2(new_n776), .B1(new_n768), .B2(new_n788), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n774), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n1054));
  INV_X1    g0854(.A(G322), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1054), .B1(new_n819), .B2(new_n784), .C1(new_n1055), .C2(new_n821), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1052), .B1(new_n600), .B2(new_n765), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n773), .A2(new_n202), .B1(new_n771), .B2(new_n246), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G150), .B2(new_n983), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n288), .B1(G97), .B2(new_n829), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n769), .A2(new_n578), .B1(new_n777), .B2(G77), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n762), .A2(new_n821), .B1(new_n819), .B2(new_n467), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1061), .A2(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n750), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n700), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n799), .A2(new_n1071), .B1(new_n254), .B2(new_n697), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n237), .A2(new_n312), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n576), .A2(G50), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT50), .Z(new_n1075));
  OAI211_X1 g0875(.A(new_n700), .B(new_n312), .C1(new_n246), .C2(new_n205), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n802), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1072), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n749), .B1(new_n1078), .B2(new_n798), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1070), .B(new_n1079), .C1(new_n693), .C2(new_n796), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1016), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n698), .B1(new_n993), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n737), .A2(new_n1016), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1080), .B1(new_n742), .B2(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(G393));
  OAI21_X1  g0884(.A(new_n798), .B1(new_n395), .B2(new_n214), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n803), .A2(new_n244), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n748), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n756), .A2(G150), .B1(G159), .B2(new_n774), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n765), .A2(new_n425), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n768), .A2(new_n205), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G68), .C2(new_n777), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n771), .A2(new_n576), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n288), .B(new_n1093), .C1(G143), .C2(new_n983), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(new_n819), .C2(new_n202), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n756), .A2(G317), .B1(G311), .B2(new_n774), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n389), .B1(new_n771), .B2(new_n832), .C1(new_n254), .C2(new_n765), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G116), .B2(new_n769), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n776), .A2(new_n788), .B1(new_n761), .B2(new_n1055), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT113), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(new_n819), .C2(new_n617), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1089), .A2(new_n1095), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1087), .B1(new_n1103), .B2(new_n750), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n997), .B2(new_n796), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1012), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n742), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n699), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  NAND2_X1  g0911(.A1(new_n922), .A2(new_n923), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n879), .A2(new_n926), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n879), .A2(new_n926), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n925), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n684), .B1(new_n939), .B2(new_n944), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n935), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n935), .B(G330), .C1(new_n727), .C2(new_n734), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1113), .B(new_n1120), .C1(new_n1114), .C2(new_n925), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n743), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n749), .B1(new_n467), .B2(new_n811), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n756), .A2(G128), .B1(G132), .B2(new_n774), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT115), .Z(new_n1127));
  NOR2_X1   g0927(.A1(new_n776), .A2(new_n468), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n768), .A2(new_n762), .B1(new_n765), .B2(new_n202), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n268), .B1(new_n761), .B2(new_n1131), .C1(new_n771), .C2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1130), .B(new_n1133), .C1(new_n757), .C2(G137), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n389), .B1(new_n776), .B2(new_n425), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT117), .Z(new_n1140));
  AOI22_X1  g0940(.A1(new_n774), .A2(G116), .B1(new_n817), .B2(G97), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n832), .B2(new_n761), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1091), .B(new_n1142), .C1(G68), .C2(new_n829), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n757), .A2(G107), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n756), .A2(G283), .ZN(new_n1145));
  AND4_X1   g0945(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1137), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1125), .B1(new_n751), .B2(new_n1147), .C1(new_n925), .C2(new_n794), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1116), .A2(new_n599), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n660), .B(new_n1151), .C1(new_n867), .C2(new_n871), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT114), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n878), .B1(new_n1116), .B2(new_n816), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n852), .A2(new_n813), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1120), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1153), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n934), .A2(G330), .A3(new_n816), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n877), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(KEYINPUT114), .A3(new_n1155), .A4(new_n1120), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n877), .B1(new_n735), .B2(new_n849), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1117), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1155), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1152), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n699), .B1(new_n1167), .B2(new_n1122), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1123), .A2(new_n1166), .A3(new_n1152), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1149), .A2(new_n1170), .ZN(G378));
  AOI21_X1  g0971(.A(new_n684), .B1(new_n945), .B2(new_n946), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n475), .A2(new_n670), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n491), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n486), .A2(new_n490), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1175), .B1(new_n486), .B2(new_n490), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n490), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1173), .B(new_n1181), .C1(new_n482), .C2(new_n485), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT120), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1178), .A2(new_n1183), .A3(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1172), .A2(new_n937), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1172), .A2(new_n937), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1184), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n929), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n903), .A2(KEYINPUT102), .B1(new_n925), .B2(new_n927), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1172), .A2(new_n937), .A3(new_n1188), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1184), .B1(new_n1172), .B2(new_n937), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n906), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT121), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1193), .A2(new_n1197), .A3(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1157), .A2(new_n1160), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1152), .B1(new_n1122), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1197), .A4(new_n1193), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n698), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G97), .A2(new_n757), .B1(new_n756), .B2(G116), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n765), .A2(new_n537), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1210), .B(new_n975), .C1(G77), .C2(new_n777), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n771), .A2(new_n437), .B1(new_n761), .B2(new_n788), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n288), .A2(new_n305), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G107), .C2(new_n774), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT119), .Z(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n776), .A2(new_n1132), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n773), .A2(new_n1220), .B1(new_n771), .B2(new_n820), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G150), .C2(new_n769), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n819), .B2(new_n827), .C1(new_n1131), .C2(new_n821), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n829), .A2(G159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n983), .C2(G124), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1213), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT118), .Z(new_n1230));
  NAND4_X1  g1030(.A1(new_n1217), .A2(new_n1218), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n750), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n745), .B1(new_n202), .B2(new_n811), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n1188), .C2(new_n794), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1202), .B2(new_n743), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1208), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n872), .A2(new_n1150), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1203), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1019), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1167), .A3(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT122), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n877), .A2(new_n793), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n750), .A2(G68), .A3(new_n793), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n773), .A2(new_n820), .B1(new_n771), .B2(new_n468), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G128), .B2(new_n983), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1210), .A2(new_n288), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n769), .A2(G50), .B1(new_n777), .B2(G159), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n827), .A2(new_n821), .B1(new_n819), .B2(new_n1132), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n600), .A2(new_n819), .B1(new_n821), .B2(new_n832), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n974), .B1(new_n578), .B2(new_n769), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n268), .B1(new_n774), .B2(G283), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G107), .A2(new_n817), .B1(new_n983), .B2(G303), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n777), .A2(G97), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1249), .A2(new_n1250), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n749), .B(new_n1244), .C1(new_n1257), .C2(new_n750), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1166), .A2(new_n743), .B1(new_n1243), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1242), .A2(new_n1259), .ZN(G381));
  OAI21_X1  g1060(.A(new_n1041), .B1(new_n1048), .B2(new_n743), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT111), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1049), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n992), .A3(new_n1110), .A4(new_n1265), .ZN(new_n1266));
  OR3_X1    g1066(.A1(G381), .A2(new_n1266), .A3(KEYINPUT123), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT123), .B1(G381), .B2(new_n1266), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1208), .A2(new_n1270), .A3(new_n1236), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1267), .A2(new_n1268), .A3(new_n1272), .ZN(G407));
  NAND3_X1  g1073(.A1(new_n673), .A2(new_n674), .A3(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(KEYINPUT124), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(KEYINPUT124), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(G213), .A3(G407), .A4(new_n1278), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1152), .B2(new_n1166), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n699), .B1(new_n1152), .B2(new_n1166), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1238), .A2(new_n1203), .A3(KEYINPUT60), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1284), .A2(G384), .A3(new_n1259), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1284), .B2(new_n1259), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G378), .B(new_n1236), .C1(new_n1205), .C2(new_n1207), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1193), .A2(new_n1197), .A3(KEYINPUT121), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT121), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1240), .B(new_n1204), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1193), .A2(new_n1197), .A3(new_n743), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1234), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1270), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1293), .B2(new_n1270), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1274), .B(new_n1287), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1297), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1288), .A3(new_n1295), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1274), .A4(new_n1287), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(new_n809), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n992), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1307), .B(new_n1110), .C1(new_n1263), .C2(new_n1049), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G390), .B1(new_n1264), .B2(new_n992), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1306), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G387), .A2(new_n1110), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1264), .A2(new_n992), .A3(G390), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1305), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1274), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1285), .A2(new_n1286), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1275), .A2(G2897), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1320), .B(new_n1323), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1321), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1318), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1316), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT127), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1302), .A2(new_n1334), .A3(new_n1274), .A4(new_n1287), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1314), .B1(new_n1332), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1331), .A2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(G375), .A2(G378), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1271), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1287), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1339), .B(new_n1271), .C1(new_n1286), .C2(new_n1285), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1315), .ZN(G402));
endmodule


