//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT74), .B1(new_n187), .B2(G104), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT74), .ZN(new_n193));
  OAI21_X1  g007(.A(G101), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n187), .A2(KEYINPUT3), .A3(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT3), .B1(new_n187), .B2(G104), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n192), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(KEYINPUT1), .A3(G146), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n199), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n198), .A3(new_n194), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(G137), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n221), .A3(new_n224), .A4(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(KEYINPUT12), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT12), .B1(new_n215), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n234), .B(KEYINPUT12), .C1(new_n215), .C2(new_n231), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n227), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n204), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n201), .B2(new_n203), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT64), .A3(new_n242), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n204), .B2(new_n242), .ZN(new_n251));
  INV_X1    g065(.A(new_n242), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n247), .A2(new_n249), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n238), .A2(KEYINPUT73), .A3(new_n198), .A4(KEYINPUT4), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n241), .A2(new_n254), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n231), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n214), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n214), .A2(new_n259), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n236), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT77), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n236), .B(KEYINPUT77), .C1(new_n264), .C2(new_n265), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n231), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n272), .B(new_n277), .C1(new_n264), .C2(new_n265), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(G469), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n236), .B(new_n272), .C1(new_n264), .C2(new_n265), .ZN(new_n280));
  INV_X1    g094(.A(new_n277), .ZN(new_n281));
  INV_X1    g095(.A(new_n265), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n262), .A2(new_n263), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  INV_X1    g100(.A(G469), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(new_n286), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(G469), .A2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n279), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G221), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n286), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G952), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(G234), .A2(G237), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT21), .B(G898), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(G902), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT87), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G214), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n200), .A2(KEYINPUT83), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT18), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(new_n224), .ZN(new_n315));
  NAND2_X1  g129(.A1(G125), .A2(G140), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G125), .A2(G140), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT72), .B1(new_n323), .B2(new_n316), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n202), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n317), .A2(new_n318), .A3(new_n202), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n313), .A2(new_n314), .A3(new_n224), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT19), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n320), .B2(new_n324), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n317), .A2(new_n318), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n202), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n322), .A3(G125), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n333), .B2(new_n339), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n341), .A2(new_n202), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n332), .A2(KEYINPUT84), .A3(new_n202), .A4(new_n334), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n337), .A2(new_n338), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n313), .B(new_n224), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n330), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G113), .B(G122), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT86), .B(G104), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n308), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n313), .A2(new_n224), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n345), .B2(KEYINPUT17), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n341), .B(new_n202), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n330), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(new_n345), .A3(new_n344), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(new_n352), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT87), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G475), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n286), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(G128), .B(G143), .Z(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G134), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT88), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n374), .B(new_n187), .C1(G116), .C2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(G116), .ZN(new_n378));
  OAI21_X1  g192(.A(G107), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n371), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n200), .A3(G128), .ZN(new_n382));
  OAI211_X1 g196(.A(G134), .B(new_n382), .C1(new_n370), .C2(new_n381), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT89), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT91), .Z(new_n391));
  OAI21_X1  g205(.A(KEYINPUT90), .B1(new_n378), .B2(new_n389), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n378), .A2(KEYINPUT90), .A3(new_n389), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n374), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G107), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n370), .A2(G134), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n395), .B(new_n376), .C1(new_n371), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n294), .A2(G217), .A3(new_n310), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n388), .B2(new_n397), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n286), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n403), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n360), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n286), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G475), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n365), .A2(KEYINPUT20), .A3(new_n366), .A4(new_n286), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n369), .A2(new_n407), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n297), .A2(new_n307), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G119), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G128), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(KEYINPUT71), .B2(KEYINPUT23), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n416), .A2(KEYINPUT71), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n205), .A2(G119), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G110), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n416), .A2(new_n419), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT24), .B(G110), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n357), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n422), .A2(G110), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n325), .A3(new_n342), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT22), .B(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n286), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n437), .A2(KEYINPUT25), .ZN(new_n438));
  INV_X1    g252(.A(G217), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(G234), .B2(new_n286), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(KEYINPUT25), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n437), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT32), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n251), .A2(new_n253), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT64), .B1(new_n248), .B2(new_n242), .ZN(new_n447));
  NOR4_X1   g261(.A1(new_n207), .A2(new_n246), .A3(new_n252), .A4(new_n243), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n226), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n219), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n217), .A2(G137), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n213), .A2(new_n225), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT2), .B(G113), .Z(new_n455));
  XNOR2_X1  g269(.A(G116), .B(G119), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(KEYINPUT66), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n455), .ZN(new_n462));
  INV_X1    g276(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n230), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT67), .B1(new_n223), .B2(new_n225), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n254), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n459), .A2(new_n460), .B1(new_n463), .B2(new_n462), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n453), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n449), .B2(new_n453), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  OAI211_X1 g288(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT28), .ZN(new_n476));
  INV_X1    g290(.A(new_n453), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n231), .B2(new_n254), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n478), .A2(new_n470), .B1(new_n473), .B2(KEYINPUT68), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT28), .B1(new_n478), .B2(new_n470), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n475), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n309), .A2(new_n310), .A3(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n195), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n453), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n454), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n493), .A3(new_n465), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n471), .A3(new_n489), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT31), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(KEYINPUT31), .A3(new_n471), .A4(new_n489), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n485), .A2(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(G472), .A2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n445), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT28), .B1(new_n472), .B2(new_n474), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n483), .B2(new_n482), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n489), .B1(new_n504), .B2(new_n475), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n497), .A2(new_n498), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT32), .B(new_n500), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(KEYINPUT70), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(new_n445), .C1(new_n499), .C2(new_n501), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G472), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n494), .A2(new_n471), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n490), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n513), .B(new_n515), .C1(new_n485), .C2(new_n490), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n478), .B(new_n470), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n482), .B1(new_n517), .B2(KEYINPUT28), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n490), .A2(new_n513), .ZN(new_n519));
  AOI21_X1  g333(.A(G902), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n512), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n444), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G214), .B1(G237), .B2(G902), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n241), .A2(new_n256), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT79), .A3(new_n255), .A4(new_n465), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g342(.A(G113), .B1(new_n463), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n415), .A3(G116), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT80), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n461), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n532), .A2(new_n199), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n241), .A2(new_n465), .A3(new_n255), .A4(new_n256), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n527), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT81), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n527), .A2(new_n533), .A3(new_n541), .A4(new_n536), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n544), .A3(new_n539), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n540), .A2(new_n546), .A3(KEYINPUT6), .A4(new_n542), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n254), .A2(G125), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(G125), .B2(new_n211), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n310), .A2(G224), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n551), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n532), .B(new_n199), .Z(new_n557));
  XNOR2_X1  g371(.A(new_n539), .B(KEYINPUT8), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n542), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n286), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G210), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n554), .A2(new_n286), .A3(new_n561), .A4(new_n559), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n525), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n414), .A2(new_n523), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT92), .B(G101), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(G3));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n369), .A2(new_n411), .A3(new_n412), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT33), .B1(new_n401), .B2(new_n402), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n388), .A2(new_n397), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n398), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n400), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(G478), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(G478), .A2(G902), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n404), .B(new_n286), .C1(new_n401), .C2(new_n402), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n307), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n565), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n569), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT93), .B1(new_n570), .B2(new_n579), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n307), .B(new_n525), .C1(new_n563), .C2(new_n564), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT94), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n286), .B1(new_n505), .B2(new_n506), .ZN(new_n594));
  INV_X1    g408(.A(new_n499), .ZN(new_n595));
  AOI22_X1  g409(.A1(G472), .A2(new_n594), .B1(new_n595), .B2(new_n500), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n444), .A2(new_n295), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n292), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NAND2_X1  g415(.A1(new_n563), .A2(new_n564), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n403), .B(new_n405), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n603), .A2(new_n369), .A3(new_n411), .A4(new_n412), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n602), .A2(new_n585), .A3(new_n524), .A4(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n565), .A2(KEYINPUT95), .A3(new_n585), .A4(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n598), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n430), .B(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n614), .B(new_n286), .C1(new_n439), .C2(G234), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n442), .A2(KEYINPUT96), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT96), .B1(new_n442), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n525), .B(new_n618), .C1(new_n563), .C2(new_n564), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n414), .A3(new_n596), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT37), .B(G110), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G12));
  AOI21_X1  g436(.A(new_n521), .B1(new_n508), .B2(new_n510), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n297), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n369), .A2(new_n603), .A3(new_n411), .A4(new_n412), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n301), .B1(new_n305), .B2(G900), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n205), .ZN(G30));
  NAND3_X1  g446(.A1(new_n570), .A2(new_n603), .A3(new_n524), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n442), .A2(new_n615), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n514), .A2(new_n489), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n286), .B1(new_n517), .B2(new_n489), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n511), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n297), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n627), .B(KEYINPUT39), .Z(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n602), .B(KEYINPUT38), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n643), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G143), .ZN(G45));
  NAND3_X1  g467(.A1(new_n570), .A2(new_n579), .A3(new_n627), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n625), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n202), .ZN(G48));
  NAND2_X1  g470(.A1(new_n285), .A2(new_n286), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G469), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n296), .A3(new_n290), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n523), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n584), .A2(new_n586), .A3(new_n569), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT94), .B1(new_n590), .B2(new_n591), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT98), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n593), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n669), .B(new_n671), .ZN(G15));
  AOI21_X1  g486(.A(new_n661), .B1(new_n607), .B2(new_n608), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n373), .ZN(G18));
  AOI21_X1  g488(.A(new_n413), .B1(new_n511), .B2(new_n522), .ZN(new_n675));
  INV_X1    g489(.A(new_n618), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n659), .A2(new_n307), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n565), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  OR2_X1    g493(.A1(new_n518), .A2(new_n489), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n497), .A2(new_n498), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n501), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n594), .A2(G472), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n594), .A2(new_n685), .A3(G472), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n444), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n677), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n563), .A2(new_n564), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT101), .B1(new_n690), .B2(new_n633), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n634), .A2(new_n692), .A3(new_n602), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n375), .ZN(G24));
  AOI211_X1 g509(.A(new_n635), .B(new_n682), .C1(new_n684), .C2(new_n686), .ZN(new_n696));
  INV_X1    g510(.A(new_n654), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n565), .A4(new_n660), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n563), .A2(new_n524), .A3(new_n564), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n291), .B(KEYINPUT102), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n279), .A2(new_n290), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n296), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n523), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n700), .B1(new_n707), .B2(new_n654), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n563), .A2(new_n524), .A3(new_n564), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n654), .A3(new_n705), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n502), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(KEYINPUT103), .B(new_n445), .C1(new_n499), .C2(new_n501), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n522), .A3(new_n507), .A4(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n688), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n710), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NOR4_X1   g533(.A1(new_n709), .A2(new_n623), .A3(new_n705), .A4(new_n444), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n629), .A2(KEYINPUT105), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n604), .A2(KEYINPUT105), .A3(new_n627), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n721), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n523), .A2(new_n724), .A3(new_n701), .A4(new_n706), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n726), .B2(new_n722), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  NAND4_X1  g543(.A1(new_n579), .A2(new_n411), .A3(new_n369), .A4(new_n412), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n596), .A2(new_n635), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n275), .A2(new_n278), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n275), .A2(KEYINPUT45), .A3(new_n278), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n702), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n751), .A3(KEYINPUT46), .A4(new_n703), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n747), .A2(new_n750), .A3(new_n290), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n296), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n645), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n738), .A2(new_n739), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n740), .A2(new_n701), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  XNOR2_X1  g572(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n753), .A2(new_n296), .A3(new_n759), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n709), .A2(new_n654), .A3(new_n688), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n623), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n687), .A2(new_n688), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n302), .B1(new_n732), .B2(new_n733), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n660), .B(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n650), .A2(new_n524), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n768), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n734), .A2(new_n778), .A3(new_n302), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(KEYINPUT50), .A3(new_n660), .A4(new_n775), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n709), .A2(new_n659), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n696), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n444), .A2(new_n301), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n642), .A3(new_n787), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n788), .A2(new_n570), .A3(new_n579), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n770), .A3(new_n701), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n781), .A2(new_n793), .A3(new_n701), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n658), .A2(new_n290), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(new_n296), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n761), .A2(new_n762), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n767), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n565), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT118), .B1(new_n774), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n781), .A2(new_n804), .A3(new_n565), .A4(new_n660), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n299), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n714), .A2(new_n688), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n784), .A2(new_n808), .A3(new_n785), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT119), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n784), .A2(new_n811), .A3(new_n808), .A4(new_n785), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n810), .A2(KEYINPUT48), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n807), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n799), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n792), .A2(new_n794), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n799), .A2(new_n817), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n783), .A2(new_n786), .A3(new_n789), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n825), .A4(KEYINPUT51), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n816), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n788), .A2(new_n584), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n580), .A2(new_n626), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n598), .A3(new_n565), .A4(new_n585), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n620), .A2(new_n566), .A3(new_n678), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n673), .A3(new_n694), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n667), .B1(new_n593), .B2(new_n662), .ZN(new_n833));
  AOI211_X1 g647(.A(KEYINPUT98), .B(new_n661), .C1(new_n587), .C2(new_n592), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n696), .A2(new_n697), .A3(new_n706), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n624), .A2(new_n676), .A3(new_n627), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(new_n413), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n701), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n718), .A2(new_n728), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT112), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n718), .A2(new_n728), .A3(new_n839), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n669), .A3(new_n843), .A4(new_n832), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n619), .B(new_n624), .C1(new_n629), .C2(new_n697), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(new_n698), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n691), .A2(new_n693), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n642), .A2(new_n705), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n635), .A3(new_n627), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT113), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT113), .B1(new_n848), .B2(new_n851), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n851), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT113), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT53), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n845), .A2(new_n863), .A3(new_n854), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n835), .A2(new_n840), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n854), .A4(new_n864), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n854), .A2(new_n859), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n841), .B2(new_n844), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n867), .B(new_n869), .C1(new_n871), .C2(KEYINPUT53), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n827), .A2(new_n828), .A3(new_n866), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n298), .A2(new_n310), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT110), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n597), .A2(new_n524), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n730), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n642), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n650), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n881), .B(new_n883), .C1(new_n878), .C2(new_n879), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n884), .ZN(G75));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n845), .B2(new_n860), .ZN(new_n886));
  INV_X1    g700(.A(new_n869), .ZN(new_n887));
  OAI211_X1 g701(.A(G210), .B(G902), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n548), .A2(new_n549), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n553), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n890), .B(new_n891), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n310), .A2(G952), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT123), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n869), .B1(new_n871), .B2(KEYINPUT53), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(KEYINPUT121), .A3(G210), .A4(G902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n899), .B1(new_n904), .B2(new_n892), .ZN(G51));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n886), .B2(new_n887), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n872), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n702), .B(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n285), .ZN(new_n910));
  OAI211_X1 g724(.A(G902), .B(new_n749), .C1(new_n886), .C2(new_n887), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n896), .B1(new_n910), .B2(new_n913), .ZN(G54));
  NOR2_X1   g728(.A1(new_n886), .A2(new_n887), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n286), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(new_n365), .ZN(new_n917));
  INV_X1    g731(.A(new_n896), .ZN(new_n918));
  INV_X1    g732(.A(new_n365), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n902), .A2(KEYINPUT58), .A3(G902), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n366), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(G60));
  NAND2_X1  g736(.A1(new_n571), .A2(new_n575), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n866), .A2(new_n872), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n577), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n906), .B2(new_n872), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n897), .A3(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n902), .A2(new_n932), .B1(new_n435), .B2(new_n436), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n902), .A2(new_n614), .A3(new_n932), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n898), .A4(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n898), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n310), .B1(new_n303), .B2(G224), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n835), .B2(new_n310), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT125), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n889), .B1(G898), .B2(new_n310), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AND2_X1   g759(.A1(new_n757), .A2(new_n765), .ZN(new_n946));
  INV_X1    g760(.A(new_n647), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(new_n523), .A3(new_n701), .A4(new_n829), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n652), .A2(new_n848), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n946), .A2(KEYINPUT127), .A3(new_n948), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n491), .A2(new_n493), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n332), .A2(new_n334), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT126), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n310), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(G900), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n960), .B2(new_n270), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n718), .A2(new_n728), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n755), .A2(new_n849), .A3(new_n808), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n946), .A2(new_n964), .A3(new_n848), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n310), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(G227), .B2(new_n310), .ZN(new_n968));
  OAI221_X1 g782(.A(new_n961), .B1(new_n310), .B2(new_n963), .C1(new_n960), .C2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n956), .B2(new_n835), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n639), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n966), .B2(new_n835), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n514), .A2(new_n489), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n896), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n862), .A2(new_n865), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n977), .A2(new_n638), .A3(new_n971), .A4(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n973), .A2(new_n976), .A3(new_n979), .ZN(G57));
endmodule


