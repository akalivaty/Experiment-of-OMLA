//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G197gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT11), .B(G169gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT12), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G15gat), .B(G22gat), .Z(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G1gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n215), .A3(KEYINPUT96), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT97), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT92), .B(G29gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G36gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT91), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n222), .B(new_n224), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n221), .B(new_n225), .C1(new_n226), .C2(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT15), .B1(new_n228), .B2(G43gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(G43gat), .B2(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n228), .A2(G43gat), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT93), .B(G43gat), .Z(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G50gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT15), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n226), .A2(new_n221), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n236), .A2(KEYINPUT94), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT94), .B1(new_n236), .B2(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT95), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT95), .B(new_n231), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n219), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n248), .B2(new_n218), .ZN(new_n249));
  NAND2_X1  g048(.A1(G229gat), .A2(G233gat), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT18), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n218), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n246), .B2(new_n247), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  INV_X1    g053(.A(new_n250), .ZN(new_n255));
  NOR4_X1   g054(.A1(new_n253), .A2(new_n254), .A3(new_n244), .A4(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n250), .B(KEYINPUT13), .ZN(new_n258));
  INV_X1    g057(.A(new_n244), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n242), .A2(new_n243), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n219), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n209), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NOR4_X1   g063(.A1(new_n251), .A2(new_n256), .A3(new_n262), .A4(new_n208), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n250), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  INV_X1    g067(.A(new_n256), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n263), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n208), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n263), .A3(new_n209), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(KEYINPUT98), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G228gat), .A2(G233gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G197gat), .B(G204gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT22), .ZN(new_n277));
  INV_X1    g076(.A(G211gat), .ZN(new_n278));
  INV_X1    g077(.A(G218gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G211gat), .B(G218gat), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT73), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT2), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(G148gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(G141gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT79), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n291), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300));
  INV_X1    g099(.A(new_n291), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n286), .B2(G141gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n288), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n294), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n291), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n292), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n304), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n309), .A2(new_n292), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n310), .A2(new_n317), .B1(new_n296), .B2(new_n303), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n283), .A2(new_n313), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n305), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n275), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n311), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n319), .A2(KEYINPUT85), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n305), .B1(new_n319), .B2(KEYINPUT85), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(G228gat), .A3(G233gat), .A4(new_n315), .ZN(new_n326));
  INV_X1    g125(.A(G22gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n321), .B2(new_n326), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT31), .B(G50gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(KEYINPUT86), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n328), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n328), .A2(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT71), .B(G71gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT64), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT67), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G127gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(G134gat), .ZN(new_n351));
  INV_X1    g150(.A(G134gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n351), .B(new_n353), .C1(KEYINPUT1), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT68), .ZN(new_n356));
  INV_X1    g155(.A(G120gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G113gat), .ZN(new_n358));
  INV_X1    g157(.A(G113gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G120gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n353), .A4(new_n351), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n361), .A2(new_n367), .A3(new_n362), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT69), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n361), .A2(new_n367), .A3(new_n370), .A4(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n374));
  AND2_X1   g173(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT27), .B(G183gat), .Z(new_n381));
  OAI21_X1  g180(.A(KEYINPUT28), .B1(new_n381), .B2(G190gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n389));
  OR3_X1    g188(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n380), .A2(new_n382), .A3(new_n383), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT66), .B(G183gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400));
  INV_X1    g199(.A(G169gat), .ZN(new_n401));
  INV_X1    g200(.A(G176gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n388), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT25), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n404), .A2(new_n403), .B1(new_n386), .B2(new_n387), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  INV_X1    g208(.A(G183gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n397), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n373), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n397), .B1(new_n375), .B2(new_n376), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n394), .A3(new_n395), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n409), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  AND4_X1   g217(.A1(new_n409), .A2(new_n412), .A3(new_n388), .A4(new_n405), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(new_n392), .B1(new_n366), .B2(new_n372), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n346), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n344), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  INV_X1    g224(.A(new_n346), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n373), .A2(new_n414), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n356), .A2(new_n365), .B1(new_n369), .B2(new_n371), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n392), .A3(new_n420), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n422), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n424), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT72), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n424), .A2(new_n433), .A3(new_n432), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n430), .A2(new_n431), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n344), .A2(new_n423), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n415), .A2(new_n421), .A3(new_n346), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n340), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n414), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n454), .B(KEYINPUT74), .Z(new_n455));
  NAND3_X1  g254(.A1(new_n420), .A2(KEYINPUT75), .A3(new_n392), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(KEYINPUT29), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n414), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n284), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n456), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT75), .B1(new_n420), .B2(new_n392), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n420), .A2(new_n455), .A3(new_n392), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n284), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT76), .B(G8gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(G36gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n462), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n462), .A2(new_n467), .A3(KEYINPUT30), .A4(new_n472), .ZN(new_n478));
  INV_X1    g277(.A(new_n458), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n453), .B2(new_n456), .ZN(new_n480));
  INV_X1    g279(.A(new_n466), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n480), .A2(new_n461), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n284), .B1(new_n457), .B2(new_n459), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n471), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n473), .A2(KEYINPUT77), .A3(new_n474), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n477), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n318), .A2(new_n366), .A3(new_n372), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n428), .A2(new_n492), .A3(new_n318), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n373), .A3(new_n312), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n428), .B2(new_n318), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n494), .A2(new_n495), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n373), .A2(new_n322), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n489), .ZN(new_n502));
  INV_X1    g301(.A(new_n495), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(KEYINPUT5), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n497), .A2(new_n507), .A3(new_n495), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n490), .A2(KEYINPUT82), .A3(new_n493), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  AND4_X1   g309(.A1(new_n492), .A2(new_n318), .A3(new_n366), .A4(new_n372), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n498), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n506), .B(new_n508), .C1(new_n509), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n509), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n497), .A2(new_n507), .A3(new_n495), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT83), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G1gat), .B(G29gat), .ZN(new_n518));
  INV_X1    g317(.A(G85gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT0), .B(G57gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(KEYINPUT6), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n524), .B(new_n505), .C1(new_n513), .C2(new_n516), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n522), .B(KEYINPUT87), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n511), .A2(new_n498), .A3(new_n510), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT82), .B1(new_n490), .B2(new_n493), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n515), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n506), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT83), .A3(new_n515), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n528), .B1(new_n534), .B2(new_n505), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n523), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n450), .A2(new_n451), .A3(new_n488), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n524), .B1(new_n534), .B2(new_n505), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n523), .B1(new_n527), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n539), .A2(new_n540), .A3(new_n488), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n539), .B2(new_n488), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(new_n449), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n537), .B1(new_n543), .B2(new_n451), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n497), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT39), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n503), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n501), .A2(new_n548), .A3(new_n495), .A4(new_n489), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n549), .A2(KEYINPUT39), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT88), .B1(new_n502), .B2(new_n503), .ZN(new_n551));
  INV_X1    g350(.A(new_n497), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n512), .B2(new_n509), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n551), .C1(new_n553), .C2(new_n495), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n554), .A3(new_n528), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT40), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n547), .A2(new_n554), .A3(new_n559), .A4(new_n528), .ZN(new_n560));
  INV_X1    g359(.A(new_n528), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n517), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n487), .A2(new_n558), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT37), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n460), .A2(new_n284), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n465), .A2(new_n461), .A3(new_n466), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT37), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n564), .A2(new_n471), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n523), .B(new_n570), .C1(new_n527), .C2(new_n535), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT37), .B1(new_n482), .B2(new_n483), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n564), .A2(new_n471), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n473), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n563), .B(new_n340), .C1(new_n571), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n446), .A2(KEYINPUT36), .A3(new_n448), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n447), .B1(new_n438), .B2(new_n441), .ZN(new_n578));
  INV_X1    g377(.A(new_n441), .ZN(new_n579));
  AOI211_X1 g378(.A(new_n579), .B(new_n445), .C1(new_n435), .C2(new_n437), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n340), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n541), .B2(new_n542), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n274), .B1(new_n544), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT99), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT100), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G71gat), .B(G78gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(G57gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n604), .A3(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n600), .A2(KEYINPUT103), .A3(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  INV_X1    g411(.A(G99gat), .ZN(new_n613));
  INV_X1    g412(.A(G106gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT8), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT105), .B(G92gat), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n612), .B(new_n615), .C1(G85gat), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n600), .A2(new_n605), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n619), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g422(.A(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n606), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n592), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n591), .B1(new_n622), .B2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n590), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT109), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(KEYINPUT108), .B2(new_n628), .ZN(new_n631));
  INV_X1    g430(.A(new_n590), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n631), .B(new_n632), .C1(KEYINPUT108), .C2(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT102), .ZN(new_n636));
  XNOR2_X1  g435(.A(G127gat), .B(G155gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n219), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(G183gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n410), .A3(new_n219), .ZN(new_n643));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n278), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n642), .A2(new_n643), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n644), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(new_n646), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n639), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n646), .A3(new_n652), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n638), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  AND2_X1   g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n662), .B(new_n664), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n260), .B2(new_n624), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n619), .B1(new_n246), .B2(new_n247), .ZN(new_n668));
  XOR2_X1   g467(.A(G190gat), .B(G218gat), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n667), .B2(new_n668), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n665), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n676), .A3(new_n665), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n634), .B(new_n660), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n587), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n539), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n211), .ZN(G1324gat));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n488), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT42), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n217), .B2(new_n684), .ZN(G1325gat));
  INV_X1    g487(.A(G15gat), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n681), .A2(new_n689), .A3(new_n582), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n578), .A2(new_n580), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n587), .A2(new_n691), .A3(new_n680), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n681), .A2(new_n340), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n679), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n677), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n544), .B2(new_n586), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n539), .A2(new_n488), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT84), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n539), .A2(new_n540), .A3(new_n488), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n340), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n583), .B1(new_n706), .B2(KEYINPUT110), .ZN(new_n707));
  OAI211_X1 g506(.A(KEYINPUT110), .B(new_n584), .C1(new_n541), .C2(new_n542), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n544), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n701), .A3(new_n698), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n585), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n583), .A3(new_n708), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n699), .B1(new_n716), .B2(new_n544), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(KEYINPUT111), .A3(new_n701), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n702), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n660), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n634), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n271), .A2(new_n272), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n702), .ZN(new_n725));
  AND4_X1   g524(.A1(KEYINPUT111), .A2(new_n710), .A3(new_n701), .A4(new_n698), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n717), .B2(new_n701), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(new_n723), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n539), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n220), .ZN(new_n733));
  INV_X1    g532(.A(new_n274), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n700), .A2(new_n734), .A3(new_n721), .ZN(new_n735));
  INV_X1    g534(.A(new_n539), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n732), .A2(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI221_X1 g541(.A(KEYINPUT113), .B1(new_n738), .B2(new_n739), .C1(new_n732), .C2(new_n733), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1328gat));
  INV_X1    g543(.A(G36gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n735), .A2(new_n745), .A3(new_n487), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n488), .B1(new_n724), .B2(new_n731), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n745), .ZN(G1329gat));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n691), .A3(new_n233), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n719), .A2(new_n582), .A3(new_n723), .ZN(new_n752));
  OAI211_X1 g551(.A(KEYINPUT47), .B(new_n751), .C1(new_n752), .C2(new_n233), .ZN(new_n753));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  INV_X1    g553(.A(new_n582), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n719), .A2(KEYINPUT112), .A3(new_n723), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n233), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n760), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n228), .A3(new_n584), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n340), .B1(new_n724), .B2(new_n731), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT115), .B(new_n762), .C1(new_n763), .C2(new_n228), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n584), .B1(new_n756), .B2(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(G50gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n719), .A2(new_n340), .A3(new_n723), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT48), .B(new_n762), .C1(new_n770), .C2(new_n228), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1331gat));
  INV_X1    g571(.A(new_n722), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n710), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n634), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n774), .A2(new_n660), .A3(new_n698), .A4(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n539), .B(KEYINPUT116), .Z(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n603), .ZN(G1332gat));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n487), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT49), .B(G64gat), .Z(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n780), .B2(new_n782), .ZN(G1333gat));
  AOI21_X1  g582(.A(G71gat), .B1(new_n776), .B2(new_n691), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n776), .A2(G71gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n755), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g586(.A1(new_n776), .A2(new_n584), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n660), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n719), .A2(new_n775), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n792), .A2(new_n519), .A3(new_n539), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n717), .A2(new_n773), .A3(new_n660), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n775), .ZN(new_n799));
  AOI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n736), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n793), .A2(new_n800), .ZN(G1336gat));
  NAND2_X1  g600(.A1(new_n791), .A2(new_n487), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n616), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n775), .A2(G92gat), .A3(new_n488), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n803), .B(new_n804), .C1(new_n798), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n802), .A2(new_n616), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n804), .ZN(G1337gat));
  NOR3_X1   g611(.A1(new_n792), .A2(new_n613), .A3(new_n582), .ZN(new_n813));
  AOI21_X1  g612(.A(G99gat), .B1(new_n799), .B2(new_n691), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n791), .A2(G106gat), .A3(new_n584), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n634), .B1(new_n796), .B2(new_n797), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n614), .B1(new_n817), .B2(new_n340), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(KEYINPUT53), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT118), .B(new_n821), .C1(new_n816), .C2(new_n818), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(G1339gat));
  NAND2_X1  g622(.A1(new_n620), .A2(new_n626), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n824), .B2(new_n591), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(new_n627), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT119), .B(new_n632), .C1(new_n627), .C2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n827), .A3(new_n591), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n590), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n826), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n826), .B(KEYINPUT55), .C1(new_n828), .C2(new_n831), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n834), .A2(new_n633), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n722), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n261), .A2(new_n259), .A3(new_n258), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n249), .B2(new_n250), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n265), .B1(new_n207), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n634), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n698), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n679), .A2(new_n678), .A3(new_n840), .A4(new_n836), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n660), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n680), .A2(new_n773), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n777), .A2(new_n488), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n450), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n359), .A3(new_n722), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n449), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n539), .A2(new_n487), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n274), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n357), .A3(new_n634), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n855), .B2(new_n775), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  AND2_X1   g659(.A1(new_n348), .A2(new_n350), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n853), .A2(new_n861), .A3(new_n720), .A4(new_n854), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n850), .B2(new_n720), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n698), .A2(new_n352), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n849), .A2(KEYINPUT56), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n855), .B2(new_n699), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT56), .B1(new_n849), .B2(new_n866), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n582), .A2(new_n854), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n680), .A2(new_n773), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n266), .A2(new_n836), .A3(new_n273), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n698), .B1(new_n874), .B2(new_n841), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n660), .B1(new_n875), .B2(new_n843), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(KEYINPUT121), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(new_n660), .C1(new_n875), .C2(new_n843), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n872), .B(new_n340), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n846), .B2(new_n584), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n871), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n288), .B1(new_n884), .B2(new_n722), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n755), .A2(new_n340), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n846), .A2(new_n847), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G141gat), .A3(new_n274), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT58), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n871), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n734), .B(new_n890), .C1(new_n880), .C2(new_n882), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT58), .B1(new_n891), .B2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n888), .B(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n892), .A2(KEYINPUT123), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(new_n887), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n286), .A3(new_n634), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n680), .A2(new_n902), .A3(new_n274), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n680), .B2(new_n274), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n876), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n901), .B(new_n872), .C1(new_n906), .C2(new_n340), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n846), .A2(KEYINPUT57), .A3(new_n584), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n340), .B1(new_n905), .B2(new_n876), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT125), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n634), .A3(new_n890), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n900), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n286), .C1(new_n884), .C2(new_n634), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n899), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  AOI21_X1  g714(.A(G155gat), .B1(new_n898), .B2(new_n720), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n720), .A2(G155gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n884), .B2(new_n917), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n898), .B2(new_n698), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n698), .A2(G162gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n884), .B2(new_n920), .ZN(G1347gat));
  INV_X1    g720(.A(new_n777), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n853), .A2(new_n487), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n274), .ZN(new_n924));
  NOR4_X1   g723(.A1(new_n852), .A2(new_n736), .A3(new_n488), .A4(new_n449), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n401), .A3(new_n722), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  NOR3_X1   g726(.A1(new_n923), .A2(new_n402), .A3(new_n775), .ZN(new_n928));
  AOI21_X1  g727(.A(G176gat), .B1(new_n925), .B2(new_n634), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  INV_X1    g729(.A(new_n381), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n925), .A2(new_n931), .A3(new_n720), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n923), .A2(new_n660), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n398), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n923), .B2(new_n699), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n925), .A2(new_n397), .A3(new_n698), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n777), .A2(new_n755), .A3(new_n488), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n911), .A2(G197gat), .A3(new_n734), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n852), .A2(new_n736), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n487), .A3(new_n886), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n204), .B1(new_n943), .B2(new_n773), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n941), .A2(KEYINPUT126), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1352gat));
  XOR2_X1   g748(.A(KEYINPUT127), .B(G204gat), .Z(new_n950));
  NOR3_X1   g749(.A1(new_n943), .A2(new_n775), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n911), .A2(new_n634), .A3(new_n940), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  OR3_X1    g754(.A1(new_n943), .A2(G211gat), .A3(new_n660), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n911), .A2(new_n720), .A3(new_n940), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  NAND4_X1  g759(.A1(new_n911), .A2(G218gat), .A3(new_n698), .A4(new_n940), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n279), .B1(new_n943), .B2(new_n699), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


