//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n212), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n206), .B1(new_n210), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT74), .ZN(new_n248));
  INV_X1    g0048(.A(G200), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n207), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n252), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n255), .B1(new_n262), .B2(new_n222), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G238), .A3(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G232), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G107), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n265), .B(new_n267), .C1(new_n264), .C2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n263), .A2(KEYINPUT71), .B1(new_n273), .B2(new_n250), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n255), .B(new_n275), .C1(new_n222), .C2(new_n262), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n249), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G20), .A2(G77), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT70), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n208), .A2(KEYINPUT70), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT15), .B(G87), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n278), .B1(new_n279), .B2(new_n281), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(new_n203), .B2(new_n283), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n207), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n288), .A2(new_n292), .B1(new_n221), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n291), .A2(new_n207), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .A3(new_n289), .A4(new_n293), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n289), .A2(new_n207), .A3(new_n291), .A4(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n252), .A2(G20), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n297), .A2(new_n300), .A3(G77), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n248), .B1(new_n277), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n273), .A2(new_n250), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n276), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(new_n303), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n274), .A2(G190), .A3(new_n276), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n313), .B2(new_n307), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n274), .A2(new_n315), .A3(new_n276), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g0118(.A(new_n318), .B(KEYINPUT75), .Z(new_n319));
  INV_X1    g0119(.A(new_n298), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G50), .A3(new_n301), .ZN(new_n321));
  INV_X1    g0121(.A(new_n279), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n284), .A3(new_n285), .ZN(new_n323));
  INV_X1    g0123(.A(G50), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(new_n211), .A3(new_n212), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n292), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n321), .B1(G50), .B2(new_n293), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT9), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n262), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G226), .ZN(new_n333));
  INV_X1    g0133(.A(G223), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(G222), .B2(G1698), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n260), .B1(new_n336), .B2(new_n264), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G77), .B2(new_n264), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n338), .A3(new_n255), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G200), .B2(new_n339), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n329), .A2(new_n330), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n331), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT10), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n313), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n329), .B(new_n346), .C1(G179), .C2(new_n339), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n264), .B2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G33), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n212), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT79), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT79), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(G58), .A3(G68), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(new_n213), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(G159), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n281), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n349), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n362), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n283), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n264), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n350), .B1(new_n370), .B2(new_n208), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n352), .A2(new_n354), .A3(new_n369), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n283), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(new_n350), .A3(new_n208), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G68), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n367), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n366), .B(new_n292), .C1(new_n376), .C2(new_n349), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n279), .B1(new_n252), .B2(G20), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n320), .A2(new_n378), .B1(new_n294), .B2(new_n279), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n266), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n370), .A2(KEYINPUT80), .A3(new_n334), .A4(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  AOI21_X1  g0184(.A(G1698), .B1(new_n372), .B2(new_n373), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(G223), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n250), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n254), .B1(new_n332), .B2(G232), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n313), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n389), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n315), .B(new_n391), .C1(new_n387), .C2(new_n250), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n380), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n372), .A2(new_n373), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(G226), .A3(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n385), .A2(new_n384), .A3(G223), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(G223), .A3(new_n266), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(G190), .B(new_n389), .C1(new_n403), .C2(new_n260), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n391), .B1(new_n387), .B2(new_n250), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n249), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n395), .B1(new_n406), .B2(new_n380), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n380), .C1(new_n390), .C2(new_n392), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n377), .A2(new_n379), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n400), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n260), .B1(new_n411), .B2(new_n382), .ZN(new_n412));
  OAI21_X1  g0212(.A(G200), .B1(new_n412), .B2(new_n391), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n413), .A4(new_n404), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n394), .A2(new_n407), .A3(new_n409), .A4(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n286), .B2(new_n221), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n292), .ZN(new_n418));
  XOR2_X1   g0218(.A(new_n418), .B(KEYINPUT11), .Z(new_n419));
  NAND2_X1  g0219(.A1(new_n294), .A2(new_n212), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT12), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(new_n212), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(KEYINPUT77), .B2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n230), .A2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G226), .B2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n355), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n254), .B1(new_n431), .B2(new_n250), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n332), .A2(G238), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n432), .B2(new_n433), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n427), .B1(new_n439), .B2(G169), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n427), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n434), .A2(KEYINPUT13), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n436), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n315), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n426), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n443), .A2(new_n340), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(G200), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n425), .A4(new_n424), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR4_X1   g0249(.A1(new_n319), .A2(new_n348), .A3(new_n415), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n280), .A2(G77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT6), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n452), .A2(new_n453), .A3(G107), .ZN(new_n454));
  XNOR2_X1  g0254(.A(G97), .B(G107), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n451), .B1(new_n456), .B2(new_n208), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n351), .A2(new_n356), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n271), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT81), .B(new_n451), .C1(new_n456), .C2(new_n208), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n292), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n293), .A2(G97), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n283), .A2(G1), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n298), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT82), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT4), .B1(new_n385), .B2(G244), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n352), .A2(new_n354), .A3(G250), .A4(G1698), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT4), .A2(G244), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n352), .A2(new_n354), .A3(new_n473), .A4(new_n266), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n470), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n476), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n222), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(KEYINPUT82), .C1(new_n479), .C2(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(new_n250), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(G41), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n252), .B(G45), .C1(new_n484), .C2(KEYINPUT5), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(KEYINPUT5), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n485), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n490), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n260), .B(G257), .C1(new_n486), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n481), .A2(new_n315), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n478), .B1(new_n479), .B2(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n260), .B1(new_n497), .B2(new_n470), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(new_n480), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n469), .B(new_n496), .C1(new_n499), .C2(G169), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n481), .A2(G190), .A3(new_n495), .ZN(new_n501));
  INV_X1    g0301(.A(new_n468), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n463), .B2(new_n292), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n501), .B(new_n503), .C1(new_n499), .C2(new_n249), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n504), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT19), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n284), .A2(G97), .A3(new_n285), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n268), .A2(new_n270), .A3(new_n217), .A4(new_n453), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n208), .B1(new_n428), .B2(new_n510), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n396), .A2(new_n208), .A3(G68), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n292), .ZN(new_n517));
  INV_X1    g0317(.A(new_n287), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n293), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n298), .A2(new_n217), .A3(new_n466), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n483), .A2(new_n251), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n218), .B1(new_n482), .B2(G1), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n260), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n216), .A2(new_n266), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n222), .A2(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n370), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n250), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n249), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n509), .B1(new_n523), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n372), .B2(new_n373), .ZN(new_n536));
  INV_X1    g0336(.A(new_n528), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n250), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G190), .A3(new_n526), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n526), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n519), .B1(new_n516), .B2(new_n292), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT85), .A4(new_n522), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n535), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n224), .A2(G1698), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G257), .B2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n373), .B2(new_n372), .ZN(new_n547));
  INV_X1    g0347(.A(G303), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n264), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n250), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n260), .B(G270), .C1(new_n486), .C2(new_n492), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n491), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(KEYINPUT21), .A3(G169), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n491), .A2(new_n551), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G179), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(G33), .B2(G283), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n283), .A2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(G20), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n292), .B2(new_n560), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(G116), .B2(new_n293), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n466), .A2(new_n559), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n297), .A2(new_n300), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n552), .B(G169), .C1(new_n563), .C2(new_n565), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n556), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n467), .A2(new_n518), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n542), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n533), .A2(new_n315), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(G169), .C2(new_n533), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n552), .A2(G200), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n563), .A2(new_n565), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n340), .C2(new_n552), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n544), .A2(new_n569), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n352), .A2(new_n354), .A3(new_n208), .A4(G87), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n268), .A2(new_n270), .A3(G20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT23), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT86), .B1(new_n528), .B2(G20), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT86), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(new_n208), .A3(G33), .A4(G116), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n580), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT22), .A2(G87), .ZN(new_n589));
  AOI211_X1 g0389(.A(G20), .B(new_n589), .C1(new_n372), .C2(new_n373), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT24), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n396), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n578), .A2(new_n579), .B1(new_n581), .B2(KEYINPUT23), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n587), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n328), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n293), .A2(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  INV_X1    g0398(.A(new_n467), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n223), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n260), .B1(new_n492), .B2(new_n486), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n603), .A2(new_n224), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n396), .A2(G250), .A3(new_n266), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n396), .A2(G257), .A3(G1698), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G294), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n605), .B1(new_n609), .B2(new_n250), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n491), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n313), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n250), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(new_n315), .A3(new_n491), .A4(new_n604), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n602), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n610), .A2(new_n340), .A3(new_n491), .ZN(new_n616));
  AOI21_X1  g0416(.A(G200), .B1(new_n610), .B2(new_n491), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n577), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n450), .A2(new_n506), .A3(new_n508), .A4(new_n620), .ZN(G372));
  NAND3_X1  g0421(.A1(new_n448), .A2(new_n407), .A3(new_n414), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n317), .B2(new_n445), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n394), .A2(new_n409), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n345), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n347), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n450), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n500), .A2(new_n504), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n568), .A2(new_n567), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n567), .B(new_n313), .C1(new_n554), .C2(new_n550), .ZN(new_n631));
  INV_X1    g0431(.A(new_n555), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n566), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n614), .B1(new_n596), .B2(new_n600), .ZN(new_n634));
  AOI21_X1  g0434(.A(G169), .B1(new_n610), .B2(new_n491), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n630), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n542), .A2(new_n570), .B1(new_n533), .B2(new_n315), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n532), .B2(new_n250), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n250), .C1(new_n536), .C2(new_n537), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n526), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n313), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(G200), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n517), .A2(new_n539), .A3(new_n520), .A4(new_n522), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n637), .A2(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n629), .A2(new_n618), .A3(new_n636), .A4(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n538), .A2(KEYINPUT87), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n527), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n571), .B(new_n572), .C1(G169), .C2(new_n650), .ZN(new_n651));
  AOI211_X1 g0451(.A(new_n519), .B(new_n521), .C1(new_n516), .C2(new_n292), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n652), .B(new_n539), .C1(new_n650), .C2(new_n249), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n648), .B1(new_n500), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(G169), .B1(new_n481), .B2(new_n495), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n503), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n544), .A3(new_n496), .A4(new_n573), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n648), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n647), .A2(new_n659), .A3(new_n651), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n627), .B1(new_n628), .B2(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n252), .A2(new_n208), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G343), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT88), .Z(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n575), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n569), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT89), .B1(new_n569), .B2(new_n576), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(new_n670), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n569), .A2(KEYINPUT89), .A3(new_n576), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT90), .ZN(new_n676));
  XNOR2_X1  g0476(.A(KEYINPUT91), .B(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n669), .A2(new_n601), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n619), .A2(new_n680), .B1(new_n615), .B2(new_n669), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n633), .A2(new_n630), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n669), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n619), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n615), .A2(new_n668), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n204), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n512), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n214), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n543), .A2(new_n539), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT85), .B1(new_n652), .B2(new_n541), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n573), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n648), .B1(new_n699), .B2(new_n500), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n481), .A2(new_n315), .A3(new_n495), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n701), .A2(new_n656), .A3(new_n503), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT26), .A3(new_n646), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n634), .A2(new_n635), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n618), .B(new_n646), .C1(new_n705), .C2(new_n683), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n651), .B1(new_n706), .B2(new_n507), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n669), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n660), .B2(new_n669), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT93), .B1(new_n660), .B2(new_n669), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n709), .A2(new_n711), .B1(new_n712), .B2(KEYINPUT29), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n620), .A2(new_n506), .A3(new_n508), .A4(new_n669), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n632), .A2(new_n610), .A3(new_n533), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n481), .A2(new_n495), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n555), .A2(new_n540), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n499), .A2(KEYINPUT30), .A3(new_n610), .A4(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(G179), .B1(new_n554), .B2(new_n550), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n717), .A2(new_n611), .A3(new_n642), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n668), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n726), .A3(new_n668), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n714), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n713), .B1(new_n678), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n696), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n676), .A2(new_n678), .ZN(new_n732));
  INV_X1    g0532(.A(G13), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n252), .B1(new_n734), .B2(G45), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n732), .B(new_n679), .C1(new_n691), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n315), .A2(G200), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n208), .B1(new_n737), .B2(KEYINPUT96), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(KEYINPUT96), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G107), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n739), .A2(new_n340), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G87), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n264), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT97), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT98), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n208), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(KEYINPUT95), .B(G159), .Z(new_n751));
  NOR3_X1   g0551(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  INV_X1    g0553(.A(new_n751), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n749), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n340), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n315), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n752), .B(new_n755), .C1(G97), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G179), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n340), .A2(new_n249), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n761), .A2(new_n756), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G50), .A2(new_n763), .B1(new_n764), .B2(G58), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n340), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n249), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n761), .A2(new_n340), .A3(new_n249), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G68), .A2(new_n767), .B1(new_n769), .B2(G77), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n767), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  INV_X1    g0573(.A(new_n764), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  AOI21_X1  g0577(.A(new_n264), .B1(new_n749), .B2(G329), .ZN(new_n778));
  INV_X1    g0578(.A(new_n758), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G326), .B2(new_n763), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n769), .A2(G311), .B1(new_n740), .B2(G283), .ZN(new_n783));
  INV_X1    g0583(.A(new_n742), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n782), .B(new_n783), .C1(new_n548), .C2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n748), .A2(new_n771), .B1(new_n777), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n207), .B1(G20), .B2(new_n313), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n735), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n690), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n396), .A2(new_n689), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n214), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n482), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n243), .B2(new_n482), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n689), .A2(new_n355), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G355), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G116), .C2(new_n204), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n787), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n791), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n788), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n675), .B2(new_n802), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n736), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n668), .A2(new_n303), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n312), .A2(new_n317), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n307), .A2(new_n313), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n811), .A2(new_n668), .A3(new_n303), .A4(new_n316), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT102), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n314), .A2(new_n814), .A3(new_n316), .A4(new_n668), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n668), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n699), .A2(new_n500), .A3(new_n648), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT26), .B1(new_n702), .B2(new_n646), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n817), .B1(new_n820), .B2(new_n707), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n669), .B1(new_n820), .B2(new_n707), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n810), .A2(new_n816), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n729), .A2(new_n678), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n790), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n787), .A2(new_n800), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n790), .B1(G77), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT100), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n264), .B1(new_n749), .B2(G311), .ZN(new_n833));
  INV_X1    g0633(.A(new_n763), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n453), .B2(new_n779), .C1(new_n834), .C2(new_n548), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G294), .B2(new_n764), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n740), .A2(G87), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n767), .A2(G283), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n769), .A2(G116), .B1(new_n742), .B2(G107), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G137), .A2(new_n763), .B1(new_n764), .B2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n768), .B2(new_n751), .C1(new_n842), .C2(new_n772), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n740), .A2(G68), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n742), .A2(G50), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n758), .A2(G58), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n370), .B1(G132), .B2(new_n749), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n832), .B1(new_n851), .B2(new_n787), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n801), .B2(new_n824), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n828), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n734), .A2(new_n252), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n380), .A2(new_n666), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n415), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n410), .A2(new_n404), .A3(new_n413), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n393), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n393), .A2(new_n860), .A3(new_n863), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n376), .A2(new_n349), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n292), .B1(new_n376), .B2(new_n349), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n379), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n666), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n415), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n871), .B1(new_n390), .B2(new_n392), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n875), .A2(new_n860), .A3(new_n872), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n864), .B1(new_n876), .B2(new_n863), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n426), .A2(new_n668), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n445), .A2(new_n448), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n426), .B(new_n668), .C1(new_n440), .C2(new_n444), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n824), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n714), .B2(new_n728), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT40), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n874), .A2(new_n877), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n878), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n450), .A2(new_n729), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n677), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  INV_X1    g0698(.A(new_n883), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n317), .A2(new_n668), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n821), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n821), .A2(KEYINPUT105), .A3(new_n901), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n891), .ZN(new_n907));
  INV_X1    g0707(.A(new_n666), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n624), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n879), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n445), .A2(new_n668), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n626), .B1(new_n713), .B2(new_n450), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n916), .B(new_n917), .Z(new_n918));
  AOI21_X1  g0718(.A(new_n856), .B1(new_n898), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n898), .ZN(new_n920));
  INV_X1    g0720(.A(new_n456), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n559), .B(new_n210), .C1(new_n921), .C2(KEYINPUT35), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(KEYINPUT35), .B2(new_n921), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT36), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n794), .A2(G77), .A3(new_n361), .A4(new_n359), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n926), .A2(KEYINPUT103), .B1(new_n324), .B2(G68), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT103), .B2(new_n926), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n733), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n920), .A2(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n668), .A2(new_n523), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n651), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n646), .B2(new_n934), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n802), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n237), .A2(new_n793), .ZN(new_n939));
  INV_X1    g0739(.A(new_n803), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n689), .B2(new_n518), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n791), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n787), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n758), .A2(G68), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n774), .B2(new_n842), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G143), .B2(new_n763), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT113), .Z(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  INV_X1    g0748(.A(new_n740), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n264), .B1(new_n948), .B2(new_n750), .C1(new_n949), .C2(new_n221), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n772), .A2(new_n751), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n768), .A2(new_n324), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n784), .A2(new_n211), .ZN(new_n953));
  OR4_X1    g0753(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G303), .A2(new_n764), .B1(new_n763), .B2(G311), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT112), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n742), .A2(G116), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT46), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n370), .B1(new_n959), .B2(new_n750), .C1(new_n779), .C2(new_n272), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G97), .B2(new_n740), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G294), .A2(new_n767), .B1(new_n769), .B2(G283), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n947), .A2(new_n954), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  OAI211_X1 g0765(.A(new_n938), .B(new_n942), .C1(new_n943), .C2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n690), .B(KEYINPUT41), .Z(new_n967));
  OAI21_X1  g0767(.A(new_n629), .B1(new_n503), .B2(new_n669), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n702), .A2(new_n668), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n687), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT111), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n687), .B(new_n970), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n975), .C1(new_n970), .C2(new_n687), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n974), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n682), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n685), .ZN(new_n981));
  INV_X1    g0781(.A(new_n684), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n681), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n679), .B(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n730), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n967), .B1(new_n985), .B2(new_n730), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n789), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n682), .B1(new_n968), .B2(new_n969), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n968), .A2(new_n615), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n669), .B1(new_n989), .B2(new_n702), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT42), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n981), .B1(new_n968), .B2(new_n969), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n991), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n993), .A2(new_n994), .B1(new_n995), .B2(new_n937), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n937), .A2(new_n995), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n988), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n966), .B1(new_n987), .B2(new_n999), .ZN(G387));
  AOI22_X1  g0800(.A1(G317), .A2(new_n764), .B1(new_n763), .B2(G322), .ZN(new_n1001));
  INV_X1    g0801(.A(G311), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n548), .B2(new_n768), .C1(new_n1002), .C2(new_n772), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n742), .A2(G294), .B1(G283), .B2(new_n758), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT115), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n949), .A2(new_n559), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n396), .B(new_n1012), .C1(G326), .C2(new_n749), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n779), .A2(new_n287), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n370), .B(new_n1015), .C1(G150), .C2(new_n749), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G50), .A2(new_n764), .B1(new_n763), .B2(G159), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G77), .A2(new_n742), .B1(new_n740), .B2(G97), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n322), .A2(new_n767), .B1(new_n769), .B2(G68), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n943), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n692), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n1022), .C1(G68), .C2(G77), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n279), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n793), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n482), .B2(new_n233), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1022), .A2(new_n797), .B1(new_n223), .B2(new_n689), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT114), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n940), .B1(new_n1029), .B2(KEYINPUT114), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n791), .B(new_n1021), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT116), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n802), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n681), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n789), .B2(new_n984), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n984), .A2(new_n730), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n984), .A2(new_n730), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n690), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(G393));
  NAND2_X1  g0843(.A1(new_n980), .A2(new_n789), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n970), .A2(new_n1036), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n769), .A2(G294), .B1(new_n742), .B2(G283), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n548), .B2(new_n772), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1002), .A2(new_n774), .B1(new_n834), .B2(new_n959), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT52), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n355), .B1(new_n750), .B2(new_n775), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G116), .B2(new_n758), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n741), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n842), .A2(new_n834), .B1(new_n774), .B2(new_n364), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT51), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n779), .A2(new_n221), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n370), .B(new_n1059), .C1(G143), .C2(new_n749), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n837), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G50), .A2(new_n767), .B1(new_n769), .B2(new_n322), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n212), .B2(new_n784), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1047), .A2(new_n1054), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n787), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n803), .B1(new_n453), .B2(new_n204), .C1(new_n793), .C2(new_n246), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n790), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n985), .A2(new_n690), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n980), .B1(new_n730), .B2(new_n984), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1044), .B1(new_n1045), .B2(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(G390));
  NAND4_X1  g0870(.A1(new_n729), .A2(G330), .A3(new_n824), .A4(new_n883), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n669), .B(new_n824), .C1(new_n704), .C2(new_n707), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n901), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n883), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n913), .B1(new_n868), .B2(new_n878), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT117), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT117), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n874), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n867), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n859), .B2(new_n865), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n912), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n899), .B1(new_n1073), .B2(new_n901), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n903), .B(new_n900), .C1(new_n660), .C2(new_n817), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT105), .B1(new_n821), .B2(new_n901), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n883), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1088), .A2(new_n912), .B1(new_n911), .B2(new_n914), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1072), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n911), .A2(new_n914), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n906), .B2(new_n913), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n810), .A2(new_n816), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n677), .B(new_n1094), .C1(new_n714), .C2(new_n728), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n883), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n735), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1091), .A2(new_n800), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n355), .B1(new_n749), .B2(G125), .ZN(new_n1101));
  INV_X1    g0901(.A(G128), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1101), .B1(new_n364), .B2(new_n779), .C1(new_n834), .C2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  AOI22_X1  g0904(.A1(new_n769), .A2(new_n1104), .B1(new_n740), .B2(G50), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n948), .B2(new_n772), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(G132), .C2(new_n764), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n742), .A2(G150), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT53), .Z(new_n1109));
  AOI211_X1 g0909(.A(new_n264), .B(new_n1059), .C1(G294), .C2(new_n749), .ZN(new_n1110));
  INV_X1    g0910(.A(G283), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n834), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G116), .B2(new_n764), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n271), .A2(new_n767), .B1(new_n769), .B2(G97), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1114), .A2(new_n743), .A3(new_n845), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1107), .A2(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n790), .B1(new_n322), .B2(new_n830), .C1(new_n1116), .C2(new_n943), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT118), .Z(new_n1118));
  AOI21_X1  g0918(.A(new_n1099), .B1(new_n1100), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n904), .A2(new_n905), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1071), .B1(new_n1095), .B2(new_n883), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1074), .B1(new_n1095), .B2(new_n883), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n729), .A2(G330), .A3(new_n824), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n899), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1120), .A2(new_n1121), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n450), .A2(G330), .A3(new_n729), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT29), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n707), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n700), .A2(new_n703), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1130), .B2(new_n669), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n822), .A2(KEYINPUT93), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n822), .A2(new_n710), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1131), .A2(new_n1132), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1126), .B(new_n627), .C1(new_n1134), .C2(new_n628), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1125), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1098), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1090), .A2(new_n1097), .A3(new_n1136), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n690), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1119), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(new_n893), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n892), .B1(new_n879), .B2(new_n885), .ZN(new_n1143));
  OAI21_X1  g0943(.A(G330), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n348), .A2(new_n329), .A3(new_n666), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n329), .A2(new_n666), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n345), .A2(new_n347), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n894), .B2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n916), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n916), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n894), .A2(G330), .A3(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT121), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1135), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1139), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n1139), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n691), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT122), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT122), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1168), .B(new_n1171), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1151), .A2(new_n800), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n790), .B1(G50), .B2(new_n830), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n944), .B1(new_n834), .B2(new_n559), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT119), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n396), .A2(G41), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1111), .B2(new_n750), .C1(new_n774), .C2(new_n223), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G97), .A2(new_n767), .B1(new_n742), .B2(G77), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n740), .A2(G58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n287), .C2(new_n768), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1177), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT58), .Z(new_n1184));
  OAI22_X1  g0984(.A1(new_n774), .A2(new_n1102), .B1(new_n842), .B2(new_n779), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n769), .A2(G137), .B1(new_n742), .B2(new_n1104), .ZN(new_n1186));
  INV_X1    g0986(.A(G132), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n772), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(G125), .C2(new_n763), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n740), .A2(new_n754), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n749), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n324), .B1(G33), .B2(G41), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1184), .B1(new_n1191), .B2(new_n1195), .C1(new_n1178), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n943), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1175), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1160), .A2(new_n789), .B1(new_n1174), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1173), .A2(new_n1202), .ZN(G375));
  NAND2_X1  g1003(.A1(new_n1121), .A2(new_n1120), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n899), .A2(new_n800), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n790), .B1(G68), .B2(new_n830), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n264), .B(new_n1015), .C1(G303), .C2(new_n749), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n1111), .B2(new_n774), .C1(new_n780), .C2(new_n834), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n769), .A2(new_n271), .B1(new_n742), .B2(G97), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n221), .B2(new_n949), .C1(new_n559), .C2(new_n772), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G132), .A2(new_n763), .B1(new_n764), .B2(G137), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n370), .B1(G128), .B2(new_n749), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n324), .C2(new_n779), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n767), .A2(new_n1104), .B1(new_n742), .B2(G159), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n1181), .C1(new_n842), .C2(new_n768), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1210), .A2(new_n1212), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1208), .B1(new_n1218), .B2(new_n787), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1206), .A2(new_n789), .B1(new_n1207), .B2(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1136), .A2(new_n967), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1162), .A2(new_n1206), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  OR2_X1    g1024(.A1(G390), .A2(G384), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1224), .A2(new_n1225), .A3(G387), .A4(G381), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(G407));
  INV_X1    g1028(.A(G213), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(G343), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(new_n1231), .A3(G213), .ZN(G409));
  XNOR2_X1  g1032(.A(G393), .B(new_n807), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G387), .B(G390), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1222), .B1(new_n1137), .B2(KEYINPUT60), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1125), .A2(new_n1135), .A3(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n690), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1220), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(new_n854), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT125), .B1(new_n1245), .B2(KEYINPUT124), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1244), .B(G384), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1245), .A2(KEYINPUT124), .B1(G2897), .B2(new_n1230), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1251), .B(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1165), .A2(new_n967), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G378), .B1(new_n1254), .B2(new_n1202), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1160), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1139), .A2(new_n1162), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT121), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1139), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n690), .B1(new_n1261), .B2(KEYINPUT57), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G378), .B(new_n1202), .C1(new_n1256), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1173), .A2(KEYINPUT123), .A3(G378), .A4(new_n1202), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1255), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1253), .B1(new_n1267), .B2(new_n1230), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1267), .A2(new_n1230), .A3(new_n1245), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1240), .B(new_n1268), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1255), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1230), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1247), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1239), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1268), .A2(new_n1240), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1269), .A2(KEYINPUT63), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .A4(new_n1237), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(G405));
  XNOR2_X1  g1084(.A(new_n1237), .B(KEYINPUT126), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G375), .A2(new_n1140), .A3(new_n1119), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1272), .A2(new_n1247), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1247), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1285), .B(new_n1286), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1290), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1288), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1239), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(G402));
endmodule


