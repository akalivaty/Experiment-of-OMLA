//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT83), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT75), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G155gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT76), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n216), .B(KEYINPUT72), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n234), .A3(new_n208), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n236), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G22gat), .ZN(new_n242));
  AND2_X1   g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n243), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n207), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n205), .B(KEYINPUT83), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n244), .A2(new_n245), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G8gat), .B(G36gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G64gat), .ZN(new_n252));
  INV_X1    g051(.A(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G226gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n260), .B(new_n261), .C1(G183gat), .C2(G190gat), .ZN(new_n262));
  INV_X1    g061(.A(G169gat), .ZN(new_n263));
  INV_X1    g062(.A(G176gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n270), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  INV_X1    g073(.A(G183gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n261), .ZN(new_n281));
  INV_X1    g080(.A(new_n261), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n259), .B1(new_n282), .B2(KEYINPUT65), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n273), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n272), .B1(new_n284), .B2(new_n271), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n266), .A2(KEYINPUT26), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(new_n265), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n266), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n292));
  AOI21_X1  g091(.A(G190gat), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n276), .A3(KEYINPUT27), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT68), .B1(new_n296), .B2(KEYINPUT28), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT28), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT28), .A3(new_n277), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n285), .B1(new_n290), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n258), .B1(new_n304), .B2(KEYINPUT29), .ZN(new_n305));
  INV_X1    g104(.A(new_n272), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n282), .B1(new_n279), .B2(KEYINPUT65), .ZN(new_n307));
  INV_X1    g106(.A(new_n283), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n270), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n309), .B2(KEYINPUT25), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n298), .A2(new_n299), .ZN(new_n311));
  AOI211_X1 g110(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n293), .C2(new_n295), .ZN(new_n312));
  INV_X1    g111(.A(new_n302), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n314), .B2(new_n289), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n257), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n237), .B1(new_n305), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n257), .B1(new_n315), .B2(new_n239), .ZN(new_n318));
  INV_X1    g117(.A(new_n237), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n290), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n258), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n254), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n318), .B2(new_n321), .ZN(new_n324));
  INV_X1    g123(.A(new_n254), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n320), .B2(new_n310), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n316), .B(new_n237), .C1(new_n326), .C2(new_n257), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n328), .A2(KEYINPUT74), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT74), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n327), .A4(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n337));
  INV_X1    g136(.A(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(G127gat), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g145(.A(KEYINPUT1), .B(G127gat), .C1(new_n341), .C2(new_n343), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349));
  OAI21_X1  g148(.A(G127gat), .B1(new_n349), .B2(KEYINPUT1), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n345), .A3(new_n339), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(G134gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n348), .A2(new_n232), .A3(new_n234), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n355));
  AND3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n352), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n238), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n363), .B(KEYINPUT77), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n337), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n235), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n353), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  INV_X1    g170(.A(new_n357), .ZN(new_n372));
  INV_X1    g171(.A(new_n358), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n366), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT80), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n353), .B2(new_n355), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n368), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G1gat), .B(G29gat), .Z(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G57gat), .B(G85gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  INV_X1    g188(.A(new_n387), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n378), .A2(new_n390), .A3(new_n381), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n336), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n336), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n250), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT37), .B1(new_n317), .B2(new_n322), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT38), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT37), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n324), .A2(new_n401), .A3(new_n327), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n399), .A2(new_n400), .A3(new_n254), .A4(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n392), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n254), .A3(new_n402), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT38), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n405), .B2(KEYINPUT38), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n328), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n332), .B2(new_n335), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n365), .B1(new_n380), .B2(new_n362), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n370), .A2(new_n364), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI211_X1 g215(.A(new_n387), .B(new_n416), .C1(new_n414), .C2(new_n413), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n417), .A2(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n328), .A2(new_n329), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT74), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n328), .A2(KEYINPUT74), .A3(new_n329), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n333), .B(KEYINPUT73), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT84), .A4(new_n323), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n417), .A2(KEYINPUT40), .B1(new_n382), .B2(new_n387), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n412), .A2(new_n418), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n427), .A3(new_n249), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n315), .A2(new_n361), .ZN(new_n429));
  INV_X1    g228(.A(new_n361), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n320), .A2(new_n430), .A3(new_n310), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT64), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OR3_X1    g234(.A1(new_n432), .A2(KEYINPUT34), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n437), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT70), .B1(new_n437), .B2(KEYINPUT34), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT32), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n435), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT69), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n432), .A2(KEYINPUT69), .A3(new_n435), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n446), .ZN(new_n448));
  XNOR2_X1  g247(.A(G15gat), .B(G43gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n445), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n440), .A2(new_n446), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n440), .A2(new_n446), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n455), .B1(new_n447), .B2(new_n448), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n398), .A2(new_n428), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n336), .A2(new_n394), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n249), .A2(new_n456), .A3(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n336), .A2(new_n394), .A3(new_n395), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND4_X1   g274(.A1(new_n394), .A2(new_n249), .A3(new_n456), .A4(new_n460), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT35), .B1(new_n412), .B2(new_n425), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n475), .A2(KEYINPUT35), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT16), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(G1gat), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(G1gat), .B2(new_n480), .ZN(new_n483));
  INV_X1    g282(.A(G8gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(G71gat), .A2(G78gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(G71gat), .A2(G78gat), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n488), .A2(KEYINPUT96), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT9), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(KEYINPUT96), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n489), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n492), .B(KEYINPUT94), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n491), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n487), .A2(KEYINPUT93), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n487), .A2(KEYINPUT93), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n498), .A2(new_n486), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(KEYINPUT95), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT95), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n485), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT98), .ZN(new_n506));
  AND2_X1   g305(.A1(G231gat), .A2(G233gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G127gat), .B(G155gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT20), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n504), .ZN(new_n514));
  XOR2_X1   g313(.A(G183gat), .B(G211gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT97), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT19), .Z(new_n517));
  XOR2_X1   g316(.A(new_n514), .B(new_n517), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n512), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525));
  INV_X1    g324(.A(G85gat), .ZN(new_n526));
  AOI22_X1  g325(.A1(KEYINPUT8), .A2(new_n525), .B1(new_n526), .B2(new_n253), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n525), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n531), .A3(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(KEYINPUT100), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(KEYINPUT100), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n539), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT87), .B1(new_n548), .B2(new_n541), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT41), .ZN(new_n555));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n536), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n560));
  AND4_X1   g359(.A1(new_n559), .A2(new_n551), .A3(new_n560), .A4(new_n553), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n554), .B2(KEYINPUT17), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n551), .A2(new_n560), .A3(new_n553), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n558), .B1(new_n564), .B2(new_n535), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n277), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n556), .A2(new_n555), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT99), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G218gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n565), .A2(new_n567), .ZN(new_n574));
  OR3_X1    g373(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n569), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT90), .B1(new_n554), .B2(new_n485), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n483), .B(G8gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT90), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n580), .A2(new_n551), .A3(new_n581), .A4(new_n553), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n554), .A2(new_n485), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT13), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(KEYINPUT91), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT91), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n579), .A2(new_n582), .B1(new_n485), .B2(new_n554), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(new_n587), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n586), .B(new_n583), .C1(new_n564), .C2(new_n580), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT18), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n563), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n551), .B2(new_n553), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n597), .A2(new_n599), .A3(new_n559), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n485), .B1(new_n600), .B2(new_n561), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n601), .A2(KEYINPUT18), .A3(new_n586), .A4(new_n583), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n593), .A3(new_n602), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n603), .A2(KEYINPUT92), .A3(new_n609), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n495), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n497), .A2(new_n500), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n497), .A2(KEYINPUT95), .A3(new_n500), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT101), .B1(new_n623), .B2(new_n535), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n532), .A3(new_n530), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n503), .A2(new_n626), .A3(new_n536), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n624), .A2(new_n625), .A3(new_n632), .A4(new_n627), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n535), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(new_n264), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(G204gat), .Z(new_n638));
  OR3_X1    g437(.A1(new_n631), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n641), .B(new_n629), .C1(new_n633), .C2(new_n634), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n642), .A3(new_n631), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n638), .B(KEYINPUT102), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n479), .A2(new_n522), .A3(new_n578), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n394), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n412), .A2(new_n425), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n481), .A2(new_n484), .ZN(new_n656));
  NOR2_X1   g455(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n658), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT104), .B1(new_n658), .B2(KEYINPUT42), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(G1325gat));
  INV_X1    g461(.A(new_n469), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n649), .A2(G15gat), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(G15gat), .B1(new_n649), .B2(new_n466), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n250), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n479), .A2(new_n577), .ZN(new_n670));
  INV_X1    g469(.A(new_n522), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n648), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G29gat), .A3(new_n394), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n475), .A2(KEYINPUT35), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n476), .A2(new_n477), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n398), .A2(new_n428), .A3(new_n469), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n681), .B(new_n577), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT35), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n396), .A2(new_n397), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n473), .ZN(new_n689));
  INV_X1    g488(.A(new_n683), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n691), .B2(new_n578), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n693), .A2(new_n672), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n650), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G29gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n677), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n696), .A3(new_n697), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n673), .A2(G36gat), .A3(new_n653), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n694), .A2(new_n654), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n543), .B2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n469), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n693), .A2(new_n672), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n466), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n673), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n709), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  NAND3_X1  g515(.A1(new_n693), .A2(new_n250), .A3(new_n672), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT48), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n670), .A2(new_n204), .A3(new_n250), .A4(new_n672), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n720), .B(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n646), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n522), .A2(new_n578), .A3(new_n616), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n691), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n394), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT108), .B(G57gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n653), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n726), .A2(G71gat), .A3(new_n706), .ZN(new_n735));
  OAI21_X1  g534(.A(G71gat), .B1(new_n726), .B2(new_n469), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g537(.A1(new_n726), .A2(new_n249), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT109), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n724), .A2(G85gat), .A3(new_n394), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n616), .B1(new_n520), .B2(new_n521), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n578), .B(new_n743), .C1(new_n470), .C2(new_n478), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n578), .A4(new_n743), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n744), .A2(KEYINPUT111), .A3(new_n745), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n742), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n743), .A2(new_n646), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n693), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n394), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(G1336gat));
  OAI21_X1  g559(.A(new_n681), .B1(new_n479), .B2(new_n577), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n578), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n761), .A2(new_n654), .A3(new_n762), .A4(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT113), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n748), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n724), .A2(new_n653), .A3(G92gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n763), .A2(new_n769), .A3(G92gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n751), .A3(new_n767), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n693), .A2(new_n777), .A3(new_n654), .A4(new_n757), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(G92gat), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n775), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n776), .B1(new_n775), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n772), .B1(new_n781), .B2(new_n782), .ZN(G1337gat));
  NOR3_X1   g582(.A1(new_n706), .A2(G99gat), .A3(new_n724), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT116), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n752), .B2(new_n753), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n758), .B2(new_n469), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n693), .A2(new_n250), .A3(new_n757), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n724), .A2(G106gat), .A3(new_n249), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n749), .A2(new_n751), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n789), .A2(G106gat), .B1(new_n766), .B2(new_n793), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(new_n791), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n633), .A2(new_n629), .A3(new_n634), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n635), .B2(KEYINPUT117), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n633), .A2(new_n799), .A3(new_n629), .A4(new_n634), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT54), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n640), .B2(new_n642), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n803), .A3(new_n638), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n586), .B1(new_n601), .B2(new_n583), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n585), .A2(new_n588), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n608), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND4_X1   g608(.A1(new_n575), .A2(new_n576), .A3(new_n613), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT55), .A4(new_n638), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n806), .A2(new_n810), .A3(new_n639), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT118), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n613), .A2(new_n809), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n646), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n646), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n616), .A2(new_n639), .A3(new_n806), .A4(new_n811), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n578), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n522), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  NOR4_X1   g621(.A1(new_n522), .A2(new_n578), .A3(new_n616), .A4(new_n646), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n654), .A2(new_n394), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n473), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n617), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n616), .A2(new_n342), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT120), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n827), .B2(new_n830), .ZN(G1340gat));
  NOR2_X1   g630(.A1(new_n827), .A2(new_n724), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(new_n340), .ZN(G1341gat));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n522), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n827), .A2(new_n577), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n838));
  XOR2_X1   g637(.A(KEYINPUT56), .B(G134gat), .Z(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(G1343gat));
  INV_X1    g639(.A(G141gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n249), .B1(new_n822), .B2(new_n824), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n469), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n845), .B2(new_n617), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n812), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n646), .A2(new_n815), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n578), .B1(new_n820), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n671), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n250), .B1(new_n852), .B2(new_n823), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n842), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n854), .A2(new_n856), .A3(G141gat), .A4(new_n844), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n846), .B1(new_n857), .B2(new_n617), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1344gat));
  OR3_X1    g659(.A1(new_n845), .A2(G148gat), .A3(new_n724), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n616), .A2(new_n639), .A3(new_n806), .A4(new_n811), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n849), .A2(KEYINPUT119), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n816), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n577), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n671), .B1(new_n848), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n250), .B1(new_n867), .B2(new_n823), .ZN(new_n868));
  INV_X1    g667(.A(new_n812), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n522), .B1(new_n850), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n824), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n868), .A2(KEYINPUT57), .B1(new_n871), .B2(new_n250), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n844), .A2(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n844), .A2(KEYINPUT122), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n872), .A2(new_n646), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n856), .A3(new_n646), .A4(new_n844), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(new_n862), .A3(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n861), .B1(new_n876), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n854), .A2(new_n856), .A3(new_n844), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n222), .A3(new_n522), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n842), .A2(new_n671), .A3(new_n844), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n222), .B2(new_n882), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n880), .A2(new_n227), .A3(new_n577), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n842), .A2(new_n578), .A3(new_n844), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n227), .B2(new_n885), .ZN(G1347gat));
  AND2_X1   g685(.A1(new_n654), .A2(new_n473), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n825), .A2(new_n394), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n617), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n867), .A2(new_n823), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT123), .B1(new_n890), .B2(new_n650), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n825), .A2(new_n892), .A3(new_n394), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n263), .A3(new_n887), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n895), .B2(new_n617), .ZN(G1348gat));
  NAND4_X1  g695(.A1(new_n894), .A2(new_n264), .A3(new_n646), .A4(new_n887), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  OAI21_X1  g697(.A(G176gat), .B1(new_n888), .B2(new_n724), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  NOR2_X1   g701(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n903));
  AND2_X1   g702(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n671), .A2(new_n301), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n892), .B1(new_n825), .B2(new_n394), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT123), .B(new_n650), .C1(new_n822), .C2(new_n824), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n887), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n276), .A2(new_n278), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n888), .B2(new_n522), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n903), .B(new_n904), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  AND4_X1   g710(.A1(KEYINPUT125), .A2(new_n908), .A3(KEYINPUT60), .A4(new_n910), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1350gat));
  OR2_X1    g712(.A1(new_n888), .A2(new_n577), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n894), .A2(new_n887), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n578), .A2(new_n277), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n917), .A2(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1351gat));
  NAND2_X1  g720(.A1(new_n469), .A2(new_n654), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n249), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n891), .B2(new_n893), .ZN(new_n925));
  INV_X1    g724(.A(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n616), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n871), .A2(new_n250), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n922), .A2(new_n650), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n928), .B(new_n929), .C1(new_n842), .C2(new_n855), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n617), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n724), .A2(G204gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n872), .A2(new_n646), .A3(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G1353gat));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(new_n930), .B2(new_n522), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n872), .A2(new_n941), .A3(new_n671), .A4(new_n929), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n942), .A3(G211gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT63), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n671), .B(new_n923), .C1(new_n906), .C2(new_n907), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT126), .B1(new_n945), .B2(G211gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n925), .A2(new_n947), .A3(new_n211), .A4(new_n671), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n940), .A2(new_n942), .A3(new_n950), .A4(G211gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n949), .A3(new_n951), .ZN(G1354gat));
  NOR3_X1   g751(.A1(new_n930), .A2(new_n212), .A3(new_n577), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n925), .A2(new_n578), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n212), .ZN(G1355gat));
endmodule


