

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U552 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X2 U553 ( .A1(n752), .A2(n751), .ZN(n767) );
  OR2_X1 U554 ( .A1(n748), .A2(n722), .ZN(n725) );
  OR2_X2 U555 ( .A1(n764), .A2(n976), .ZN(n821) );
  INV_X1 U556 ( .A(KEYINPUT93), .ZN(n734) );
  NOR2_X1 U557 ( .A1(n817), .A2(KEYINPUT33), .ZN(n757) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n520) );
  OR2_X1 U559 ( .A1(n818), .A2(n817), .ZN(n518) );
  AND2_X1 U560 ( .A1(n756), .A2(n984), .ZN(n519) );
  INV_X1 U561 ( .A(KEYINPUT90), .ZN(n698) );
  XNOR2_X1 U562 ( .A(n723), .B(KEYINPUT91), .ZN(n724) );
  XNOR2_X1 U563 ( .A(n725), .B(n724), .ZN(n726) );
  INV_X1 U564 ( .A(KEYINPUT92), .ZN(n727) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n712) );
  XNOR2_X1 U566 ( .A(n713), .B(n712), .ZN(n717) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n781) );
  AND2_X2 U568 ( .A1(n525), .A2(G2104), .ZN(n870) );
  AND2_X1 U569 ( .A1(n819), .A2(n518), .ZN(n820) );
  NOR2_X1 U570 ( .A1(n633), .A2(n535), .ZN(n653) );
  XNOR2_X1 U571 ( .A(n521), .B(n520), .ZN(n869) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U573 ( .A1(n869), .A2(G137), .ZN(n524) );
  AND2_X1 U574 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  INV_X1 U576 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G101), .A2(n870), .ZN(n522) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n529) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n525), .ZN(n865) );
  NAND2_X1 U581 ( .A1(G125), .A2(n865), .ZN(n527) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n866) );
  NAND2_X1 U583 ( .A1(G113), .A2(n866), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n529), .A2(n528), .ZN(G160) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NOR2_X1 U587 ( .A1(G651), .A2(n633), .ZN(n649) );
  NAND2_X1 U588 ( .A1(G51), .A2(n649), .ZN(n532) );
  INV_X1 U589 ( .A(G651), .ZN(n535) );
  NOR2_X1 U590 ( .A1(G543), .A2(n535), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n530), .Z(n568) );
  NAND2_X1 U592 ( .A1(G63), .A2(n568), .ZN(n531) );
  NAND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U594 ( .A(KEYINPUT6), .B(n533), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n650), .A2(G89), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT4), .ZN(n537) );
  NAND2_X1 U597 ( .A1(G76), .A2(n653), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U599 ( .A(n538), .B(KEYINPUT5), .Z(n539) );
  NOR2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U601 ( .A(KEYINPUT7), .B(n541), .Z(n542) );
  XOR2_X1 U602 ( .A(KEYINPUT73), .B(n542), .Z(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(G65), .A2(n568), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT68), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G78), .A2(n653), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(n544), .Z(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U609 ( .A1(G53), .A2(n649), .ZN(n547) );
  XNOR2_X1 U610 ( .A(KEYINPUT69), .B(n547), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n650), .A2(G91), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(G299) );
  XOR2_X1 U614 ( .A(G2438), .B(G2454), .Z(n553) );
  XNOR2_X1 U615 ( .A(G2435), .B(G2430), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U617 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U618 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U620 ( .A(G2443), .B(G2446), .Z(n558) );
  XNOR2_X1 U621 ( .A(KEYINPUT100), .B(G2451), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U624 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U626 ( .A1(G68), .A2(n653), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n650), .A2(G81), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT13), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G43), .A2(n649), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n568), .A2(G56), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT71), .B(n572), .ZN(n978) );
  INV_X1 U637 ( .A(G860), .ZN(n621) );
  OR2_X1 U638 ( .A1(n978), .A2(n621), .ZN(G153) );
  INV_X1 U639 ( .A(G57), .ZN(G237) );
  INV_X1 U640 ( .A(G132), .ZN(G219) );
  INV_X1 U641 ( .A(G82), .ZN(G220) );
  NAND2_X1 U642 ( .A1(G102), .A2(n870), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n573), .B(KEYINPUT78), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n869), .A2(G138), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G126), .A2(n865), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G114), .A2(n866), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(G164) );
  NAND2_X1 U650 ( .A1(G90), .A2(n650), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G77), .A2(n653), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n582) );
  XNOR2_X1 U654 ( .A(n583), .B(n582), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G52), .A2(n649), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G64), .A2(n568), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U658 ( .A(KEYINPUT65), .B(n586), .Z(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G171) );
  NAND2_X1 U660 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n589), .B(KEYINPUT70), .ZN(n590) );
  XNOR2_X1 U662 ( .A(KEYINPUT10), .B(n590), .ZN(G223) );
  INV_X1 U663 ( .A(G223), .ZN(n833) );
  NAND2_X1 U664 ( .A1(n833), .A2(G567), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  INV_X1 U666 ( .A(G171), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G301), .A2(G868), .ZN(n592) );
  XNOR2_X1 U668 ( .A(n592), .B(KEYINPUT72), .ZN(n601) );
  INV_X1 U669 ( .A(G868), .ZN(n667) );
  NAND2_X1 U670 ( .A1(G54), .A2(n649), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G66), .A2(n568), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G92), .A2(n650), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G79), .A2(n653), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT15), .ZN(n970) );
  NAND2_X1 U678 ( .A1(n667), .A2(n970), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(G284) );
  NOR2_X1 U680 ( .A1(G286), .A2(n667), .ZN(n603) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n621), .A2(G559), .ZN(n604) );
  INV_X1 U684 ( .A(n970), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n604), .A2(n619), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(n970), .A2(n667), .ZN(n606) );
  XOR2_X1 U688 ( .A(KEYINPUT74), .B(n606), .Z(n607) );
  NOR2_X1 U689 ( .A1(G559), .A2(n607), .ZN(n609) );
  NOR2_X1 U690 ( .A1(G868), .A2(n978), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G123), .A2(n865), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n870), .A2(G99), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G135), .A2(n869), .ZN(n614) );
  NAND2_X1 U697 ( .A1(G111), .A2(n866), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n939) );
  XNOR2_X1 U700 ( .A(n939), .B(G2096), .ZN(n618) );
  INV_X1 U701 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U703 ( .A1(G559), .A2(n619), .ZN(n620) );
  XOR2_X1 U704 ( .A(n978), .B(n620), .Z(n665) );
  NAND2_X1 U705 ( .A1(n621), .A2(n665), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G55), .A2(n649), .ZN(n623) );
  NAND2_X1 U707 ( .A1(G80), .A2(n653), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G93), .A2(n650), .ZN(n624) );
  XNOR2_X1 U710 ( .A(KEYINPUT75), .B(n624), .ZN(n625) );
  NOR2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n568), .A2(G67), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n668) );
  XNOR2_X1 U714 ( .A(n629), .B(n668), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G49), .A2(n649), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U718 ( .A1(n568), .A2(n632), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G47), .A2(n649), .ZN(n637) );
  NAND2_X1 U722 ( .A1(G85), .A2(n650), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n653), .A2(G72), .ZN(n638) );
  XOR2_X1 U725 ( .A(KEYINPUT64), .B(n638), .Z(n639) );
  NOR2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n568), .A2(G60), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G88), .A2(n650), .ZN(n644) );
  NAND2_X1 U730 ( .A1(G75), .A2(n653), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G50), .A2(n649), .ZN(n646) );
  NAND2_X1 U733 ( .A1(G62), .A2(n568), .ZN(n645) );
  NAND2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n648), .A2(n647), .ZN(G166) );
  NAND2_X1 U736 ( .A1(G48), .A2(n649), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G86), .A2(n650), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U741 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n568), .A2(G61), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(G305) );
  XNOR2_X1 U744 ( .A(G288), .B(n668), .ZN(n664) );
  XOR2_X1 U745 ( .A(KEYINPUT19), .B(KEYINPUT76), .Z(n660) );
  INV_X1 U746 ( .A(G299), .ZN(n980) );
  XNOR2_X1 U747 ( .A(n980), .B(G166), .ZN(n659) );
  XNOR2_X1 U748 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U749 ( .A(n661), .B(G305), .Z(n662) );
  XNOR2_X1 U750 ( .A(G290), .B(n662), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n664), .B(n663), .ZN(n883) );
  XNOR2_X1 U752 ( .A(n665), .B(n883), .ZN(n666) );
  NOR2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n670) );
  NOR2_X1 U754 ( .A1(G868), .A2(n668), .ZN(n669) );
  NOR2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U756 ( .A(KEYINPUT77), .B(n671), .Z(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U765 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U766 ( .A1(G96), .A2(n678), .ZN(n838) );
  NAND2_X1 U767 ( .A1(n838), .A2(G2106), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U769 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U770 ( .A1(G108), .A2(n680), .ZN(n839) );
  NAND2_X1 U771 ( .A1(n839), .A2(G567), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n682), .A2(n681), .ZN(n912) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U774 ( .A1(n912), .A2(n683), .ZN(n837) );
  NAND2_X1 U775 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U776 ( .A(KEYINPUT79), .B(G166), .ZN(G303) );
  INV_X1 U777 ( .A(n781), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n780) );
  NOR2_X4 U779 ( .A1(n685), .A2(n780), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n719), .A2(G1348), .ZN(n687) );
  INV_X1 U781 ( .A(n719), .ZN(n720) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n720), .ZN(n686) );
  NOR2_X1 U783 ( .A1(n687), .A2(n686), .ZN(n692) );
  NAND2_X1 U784 ( .A1(G2072), .A2(n719), .ZN(n688) );
  XNOR2_X1 U785 ( .A(n688), .B(KEYINPUT27), .ZN(n689) );
  XNOR2_X1 U786 ( .A(KEYINPUT88), .B(n689), .ZN(n691) );
  INV_X1 U787 ( .A(G1956), .ZN(n913) );
  NOR2_X1 U788 ( .A1(n719), .A2(n913), .ZN(n690) );
  NOR2_X1 U789 ( .A1(n691), .A2(n690), .ZN(n708) );
  NAND2_X1 U790 ( .A1(n980), .A2(n708), .ZN(n702) );
  AND2_X1 U791 ( .A1(n692), .A2(n702), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n719), .A2(G1996), .ZN(n693) );
  XNOR2_X1 U793 ( .A(KEYINPUT26), .B(n693), .ZN(n697) );
  NAND2_X1 U794 ( .A1(G1341), .A2(n720), .ZN(n694) );
  XNOR2_X1 U795 ( .A(KEYINPUT89), .B(n694), .ZN(n695) );
  NOR2_X1 U796 ( .A1(n695), .A2(n978), .ZN(n696) );
  NAND2_X1 U797 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n703), .A2(n970), .ZN(n699) );
  XNOR2_X1 U799 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U800 ( .A1(n701), .A2(n700), .ZN(n707) );
  INV_X1 U801 ( .A(n702), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n703), .A2(n970), .ZN(n704) );
  AND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n980), .A2(n708), .ZN(n709) );
  XOR2_X1 U805 ( .A(n709), .B(KEYINPUT28), .Z(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n713) );
  XOR2_X1 U807 ( .A(KEYINPUT25), .B(G2078), .Z(n1006) );
  NOR2_X1 U808 ( .A1(n1006), .A2(n720), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n719), .A2(G1961), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n729) );
  OR2_X1 U811 ( .A1(n729), .A2(G301), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n746) );
  INV_X1 U813 ( .A(G8), .ZN(n718) );
  OR2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n817) );
  NOR2_X1 U815 ( .A1(G1966), .A2(n817), .ZN(n748) );
  NOR2_X1 U816 ( .A1(n720), .A2(G2084), .ZN(n744) );
  INV_X1 U817 ( .A(n744), .ZN(n721) );
  NAND2_X1 U818 ( .A1(n721), .A2(G8), .ZN(n722) );
  INV_X1 U819 ( .A(KEYINPUT30), .ZN(n723) );
  NOR2_X1 U820 ( .A1(G168), .A2(n726), .ZN(n728) );
  XNOR2_X1 U821 ( .A(n728), .B(n727), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n729), .A2(G301), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT31), .B(n732), .ZN(n745) );
  NAND2_X1 U825 ( .A1(n746), .A2(n745), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n733), .A2(G286), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n735), .B(n734), .ZN(n741) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n720), .ZN(n736) );
  XNOR2_X1 U829 ( .A(n736), .B(KEYINPUT94), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n817), .A2(G1971), .ZN(n737) );
  NOR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U832 ( .A1(G303), .A2(n739), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U835 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U836 ( .A1(G8), .A2(n744), .ZN(n750) );
  AND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n753) );
  XOR2_X1 U841 ( .A(KEYINPUT95), .B(n753), .Z(n983) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n983), .A2(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n767), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n984) );
  INV_X1 U846 ( .A(n817), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n519), .A2(n757), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n983), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n759), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U851 ( .A(KEYINPUT96), .B(n762), .Z(n764) );
  XOR2_X1 U852 ( .A(G1981), .B(KEYINPUT97), .Z(n763) );
  XNOR2_X1 U853 ( .A(G305), .B(n763), .ZN(n976) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U855 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n817), .A2(n768), .ZN(n814) );
  NAND2_X1 U858 ( .A1(G140), .A2(n869), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G104), .A2(n870), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n771), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G128), .A2(n865), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G116), .A2(n866), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U865 ( .A(KEYINPUT81), .B(n774), .ZN(n775) );
  XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n775), .ZN(n776) );
  NOR2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n779) );
  XNOR2_X1 U868 ( .A(KEYINPUT82), .B(KEYINPUT36), .ZN(n778) );
  XNOR2_X1 U869 ( .A(n779), .B(n778), .ZN(n860) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U871 ( .A1(n860), .A2(n810), .ZN(n956) );
  NOR2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n824) );
  NAND2_X1 U873 ( .A1(n956), .A2(n824), .ZN(n826) );
  INV_X1 U874 ( .A(n826), .ZN(n809) );
  NAND2_X1 U875 ( .A1(G105), .A2(n870), .ZN(n782) );
  XNOR2_X1 U876 ( .A(n782), .B(KEYINPUT38), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G141), .A2(n869), .ZN(n784) );
  NAND2_X1 U878 ( .A1(G129), .A2(n865), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G117), .A2(n866), .ZN(n785) );
  XNOR2_X1 U881 ( .A(KEYINPUT85), .B(n785), .ZN(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n849) );
  NOR2_X1 U884 ( .A1(G1996), .A2(n849), .ZN(n946) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n849), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G119), .A2(n865), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G107), .A2(n866), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U889 ( .A(KEYINPUT83), .B(n792), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G131), .A2(n869), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G95), .A2(n870), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U893 ( .A(KEYINPUT84), .B(n795), .Z(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n879) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n879), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U897 ( .A(KEYINPUT86), .B(n800), .Z(n957) );
  INV_X1 U898 ( .A(n957), .ZN(n803) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n879), .ZN(n940) );
  NOR2_X1 U901 ( .A1(n801), .A2(n940), .ZN(n802) );
  NOR2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U903 ( .A1(n946), .A2(n804), .ZN(n806) );
  XNOR2_X1 U904 ( .A(KEYINPUT39), .B(KEYINPUT98), .ZN(n805) );
  XNOR2_X1 U905 ( .A(n806), .B(n805), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n807), .A2(n824), .ZN(n808) );
  OR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n810), .A2(n860), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n811), .B(KEYINPUT99), .ZN(n959) );
  NAND2_X1 U910 ( .A1(n959), .A2(n824), .ZN(n812) );
  AND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n822) );
  AND2_X1 U912 ( .A1(n814), .A2(n822), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G1981), .A2(G305), .ZN(n815) );
  XNOR2_X1 U914 ( .A(n815), .B(KEYINPUT24), .ZN(n816) );
  XNOR2_X1 U915 ( .A(n816), .B(KEYINPUT87), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n831) );
  INV_X1 U917 ( .A(n822), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT80), .B(G1986), .Z(n823) );
  XNOR2_X1 U919 ( .A(G290), .B(n823), .ZN(n973) );
  NAND2_X1 U920 ( .A1(n957), .A2(n973), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  AND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  OR2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XOR2_X1 U926 ( .A(KEYINPUT101), .B(n834), .Z(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G188) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G325) );
  XOR2_X1 U932 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NAND2_X1 U937 ( .A1(n866), .A2(G112), .ZN(n840) );
  XOR2_X1 U938 ( .A(KEYINPUT103), .B(n840), .Z(n842) );
  NAND2_X1 U939 ( .A1(n870), .A2(G100), .ZN(n841) );
  NAND2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U941 ( .A(KEYINPUT104), .B(n843), .ZN(n848) );
  NAND2_X1 U942 ( .A1(G124), .A2(n865), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n869), .A2(G136), .ZN(n845) );
  NAND2_X1 U945 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U946 ( .A1(n848), .A2(n847), .ZN(G162) );
  XNOR2_X1 U947 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n849), .B(n939), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U950 ( .A(G160), .B(n852), .ZN(n864) );
  NAND2_X1 U951 ( .A1(G139), .A2(n869), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G103), .A2(n870), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G127), .A2(n865), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G115), .A2(n866), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n951) );
  XOR2_X1 U959 ( .A(n951), .B(G162), .Z(n862) );
  XNOR2_X1 U960 ( .A(n860), .B(G164), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n881) );
  NAND2_X1 U963 ( .A1(G130), .A2(n865), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G118), .A2(n866), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n877) );
  XNOR2_X1 U966 ( .A(KEYINPUT45), .B(KEYINPUT106), .ZN(n875) );
  NAND2_X1 U967 ( .A1(n869), .A2(G142), .ZN(n873) );
  NAND2_X1 U968 ( .A1(n870), .A2(G106), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT105), .B(n871), .Z(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U971 ( .A(n875), .B(n874), .Z(n876) );
  NOR2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U973 ( .A(n879), .B(n878), .Z(n880) );
  XNOR2_X1 U974 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U975 ( .A1(G37), .A2(n882), .ZN(G395) );
  XNOR2_X1 U976 ( .A(G286), .B(n978), .ZN(n884) );
  XNOR2_X1 U977 ( .A(n884), .B(n883), .ZN(n886) );
  XOR2_X1 U978 ( .A(n970), .B(G171), .Z(n885) );
  XNOR2_X1 U979 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U980 ( .A1(G37), .A2(n887), .ZN(G397) );
  XOR2_X1 U981 ( .A(G2100), .B(G2096), .Z(n889) );
  XNOR2_X1 U982 ( .A(KEYINPUT42), .B(G2678), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U984 ( .A(KEYINPUT43), .B(G2090), .Z(n891) );
  XNOR2_X1 U985 ( .A(G2067), .B(G2072), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U987 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U988 ( .A(G2078), .B(G2084), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(G227) );
  XOR2_X1 U990 ( .A(G1986), .B(G1971), .Z(n897) );
  XNOR2_X1 U991 ( .A(G1966), .B(G1961), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(n898), .B(G2474), .Z(n900) );
  XNOR2_X1 U994 ( .A(G1956), .B(G1981), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U996 ( .A(KEYINPUT41), .B(G1991), .Z(n902) );
  XNOR2_X1 U997 ( .A(G1996), .B(G1976), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(G229) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G397), .A2(n906), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(n912), .A2(G401), .ZN(n907) );
  XOR2_X1 U1004 ( .A(KEYINPUT107), .B(n907), .Z(n908) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(KEYINPUT108), .B(n911), .ZN(G308) );
  INV_X1 U1008 ( .A(G308), .ZN(G225) );
  INV_X1 U1009 ( .A(n912), .ZN(G319) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1011 ( .A(G20), .B(n913), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G19), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(G6), .B(G1981), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT59), .B(G4), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(KEYINPUT121), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n919), .B(G1348), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n922), .B(KEYINPUT60), .ZN(n925) );
  XOR2_X1 U1021 ( .A(G1966), .B(G21), .Z(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT122), .B(n923), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT123), .B(n926), .ZN(n928) );
  XOR2_X1 U1025 ( .A(G1961), .B(G5), .Z(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G1971), .B(G22), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G23), .B(G1976), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1030 ( .A(G1986), .B(G24), .Z(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1034 ( .A(n936), .B(KEYINPUT61), .Z(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(G16), .A2(n938), .ZN(n1026) );
  XNOR2_X1 U1037 ( .A(KEYINPUT112), .B(KEYINPUT52), .ZN(n965) );
  XOR2_X1 U1038 ( .A(G160), .B(G2084), .Z(n943) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(KEYINPUT109), .B(n941), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1042 ( .A(KEYINPUT110), .B(n944), .Z(n950) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1045 ( .A(KEYINPUT51), .B(n947), .Z(n948) );
  XNOR2_X1 U1046 ( .A(KEYINPUT111), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n962) );
  XOR2_X1 U1048 ( .A(G2072), .B(n951), .Z(n953) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1051 ( .A(KEYINPUT50), .B(n954), .Z(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT113), .B(n963), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1058 ( .A(KEYINPUT55), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n968), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .Z(n998) );
  XNOR2_X1 U1062 ( .A(G1961), .B(KEYINPUT116), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(G301), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n995) );
  XOR2_X1 U1067 ( .A(G168), .B(G1966), .Z(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n977), .Z(n993) );
  XNOR2_X1 U1070 ( .A(n978), .B(G1341), .ZN(n991) );
  XOR2_X1 U1071 ( .A(G1971), .B(G303), .Z(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT118), .B(n979), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1956), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n988) );
  INV_X1 U1075 ( .A(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT117), .B(n986), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT119), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n996), .B(KEYINPUT120), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1022) );
  XOR2_X1 U1085 ( .A(G2090), .B(G35), .Z(n1002) );
  XOR2_X1 U1086 ( .A(G2084), .B(KEYINPUT114), .Z(n999) );
  XNOR2_X1 U1087 ( .A(G34), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT54), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1015) );
  XOR2_X1 U1090 ( .A(G1991), .B(G25), .Z(n1003) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(G28), .ZN(n1012) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G33), .B(G2072), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1006), .B(G27), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1996), .B(G32), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT53), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT55), .B(n1016), .ZN(n1018) );
  INV_X1 U1103 ( .A(G29), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(G11), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT115), .B(n1020), .Z(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .Z(n1028) );
  XNOR2_X1 U1111 ( .A(KEYINPUT125), .B(n1028), .ZN(G311) );
  XOR2_X1 U1112 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

