

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737;

  OR2_X1 U372 ( .A1(n656), .A2(KEYINPUT2), .ZN(n658) );
  AND2_X1 U373 ( .A1(n396), .A2(n353), .ZN(n394) );
  AND2_X1 U374 ( .A1(n395), .A2(n573), .ZN(n353) );
  INV_X1 U375 ( .A(n512), .ZN(n554) );
  AND2_X4 U376 ( .A1(n600), .A2(n659), .ZN(n703) );
  NOR2_X2 U377 ( .A1(n643), .A2(n737), .ZN(n505) );
  XNOR2_X2 U378 ( .A(n565), .B(n564), .ZN(n734) );
  XNOR2_X2 U379 ( .A(n427), .B(n426), .ZN(n531) );
  XNOR2_X2 U380 ( .A(n493), .B(KEYINPUT35), .ZN(n609) );
  NAND2_X2 U381 ( .A1(n394), .A2(n393), .ZN(n493) );
  XNOR2_X2 U382 ( .A(n453), .B(n403), .ZN(n720) );
  XNOR2_X2 U383 ( .A(n485), .B(n401), .ZN(n453) );
  XNOR2_X1 U384 ( .A(n416), .B(n415), .ZN(n417) );
  INV_X2 U385 ( .A(G953), .ZN(n526) );
  INV_X4 U386 ( .A(G104), .ZN(n387) );
  NOR2_X1 U387 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U388 ( .A(n367), .B(n458), .ZN(n535) );
  NAND2_X2 U389 ( .A1(n370), .A2(n371), .ZN(n551) );
  XNOR2_X1 U390 ( .A(n439), .B(n438), .ZN(n602) );
  XNOR2_X1 U391 ( .A(n418), .B(n417), .ZN(n490) );
  XNOR2_X1 U392 ( .A(KEYINPUT8), .B(KEYINPUT70), .ZN(n414) );
  XNOR2_X1 U393 ( .A(n389), .B(KEYINPUT91), .ZN(n350) );
  BUF_X1 U394 ( .A(n609), .Z(n351) );
  BUF_X1 U395 ( .A(n628), .Z(n352) );
  XNOR2_X1 U396 ( .A(n389), .B(KEYINPUT91), .ZN(n515) );
  XNOR2_X2 U397 ( .A(n720), .B(G146), .ZN(n439) );
  XNOR2_X2 U398 ( .A(n368), .B(n457), .ZN(n540) );
  AND2_X2 U399 ( .A1(n531), .A2(n430), .ZN(n666) );
  XNOR2_X2 U400 ( .A(n574), .B(n548), .ZN(n677) );
  XNOR2_X1 U401 ( .A(G472), .B(KEYINPUT74), .ZN(n411) );
  NOR2_X1 U402 ( .A1(n732), .A2(n567), .ZN(n568) );
  NOR2_X1 U403 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U404 ( .A(G101), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U405 ( .A(n475), .B(n445), .ZN(n448) );
  XNOR2_X1 U406 ( .A(KEYINPUT16), .B(KEYINPUT75), .ZN(n445) );
  INV_X1 U407 ( .A(KEYINPUT82), .ZN(n455) );
  XNOR2_X1 U408 ( .A(n478), .B(n376), .ZN(n620) );
  XNOR2_X1 U409 ( .A(n479), .B(n477), .ZN(n376) );
  NAND2_X1 U410 ( .A1(n545), .A2(n662), .ZN(n358) );
  INV_X1 U411 ( .A(KEYINPUT100), .ZN(n357) );
  NOR2_X1 U412 ( .A1(n517), .A2(n494), .ZN(n573) );
  OR2_X1 U413 ( .A1(n602), .A2(n390), .ZN(n371) );
  AND2_X1 U414 ( .A1(n369), .A2(n355), .ZN(n370) );
  NAND2_X1 U415 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U416 ( .A(n512), .B(n413), .ZN(n543) );
  NAND2_X1 U417 ( .A1(n596), .A2(n595), .ZN(n600) );
  XNOR2_X1 U418 ( .A(G134), .B(G131), .ZN(n402) );
  INV_X1 U419 ( .A(KEYINPUT71), .ZN(n415) );
  XOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n522) );
  AND2_X1 U421 ( .A1(n363), .A2(n356), .ZN(n362) );
  XNOR2_X1 U422 ( .A(G902), .B(KEYINPUT15), .ZN(n593) );
  XNOR2_X1 U423 ( .A(n452), .B(n379), .ZN(n474) );
  INV_X1 U424 ( .A(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U425 ( .A(G113), .B(G143), .ZN(n477) );
  XNOR2_X1 U426 ( .A(G104), .B(G101), .ZN(n435) );
  INV_X1 U427 ( .A(KEYINPUT38), .ZN(n548) );
  INV_X1 U428 ( .A(KEYINPUT76), .ZN(n374) );
  INV_X1 U429 ( .A(G469), .ZN(n392) );
  XNOR2_X1 U430 ( .A(G134), .B(G122), .ZN(n482) );
  BUF_X1 U431 ( .A(n598), .Z(n722) );
  XNOR2_X1 U432 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT79), .ZN(n386) );
  XNOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT80), .ZN(n385) );
  XNOR2_X1 U435 ( .A(n380), .B(G125), .ZN(n452) );
  INV_X1 U436 ( .A(G146), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n451), .B(KEYINPUT81), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n449), .B(n450), .ZN(n715) );
  XNOR2_X1 U439 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U440 ( .A1(n634), .A2(n377), .ZN(n582) );
  NOR2_X1 U441 ( .A1(n378), .A2(n543), .ZN(n377) );
  INV_X1 U442 ( .A(KEYINPUT34), .ZN(n466) );
  BUF_X1 U443 ( .A(n540), .Z(n574) );
  XNOR2_X1 U444 ( .A(n375), .B(n480), .ZN(n481) );
  NOR2_X1 U445 ( .A1(n620), .A2(G902), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n425), .B(KEYINPUT25), .ZN(n426) );
  XNOR2_X1 U447 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U448 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U449 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U450 ( .A(n715), .B(n388), .ZN(n628) );
  XNOR2_X1 U451 ( .A(n383), .B(n381), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n382), .B(n452), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n453), .B(n384), .ZN(n383) );
  AND2_X1 U454 ( .A1(n605), .A2(G953), .ZN(n707) );
  XNOR2_X1 U455 ( .A(n553), .B(KEYINPUT42), .ZN(n735) );
  XNOR2_X1 U456 ( .A(n358), .B(n357), .ZN(n498) );
  NOR2_X1 U457 ( .A1(n698), .A2(G953), .ZN(n699) );
  NOR2_X1 U458 ( .A1(n695), .A2(n400), .ZN(n696) );
  AND2_X1 U459 ( .A1(n505), .A2(n507), .ZN(n354) );
  INV_X1 U460 ( .A(G902), .ZN(n391) );
  NAND2_X1 U461 ( .A1(G902), .A2(G469), .ZN(n355) );
  INV_X1 U462 ( .A(n541), .ZN(n634) );
  OR2_X1 U463 ( .A1(n507), .A2(KEYINPUT44), .ZN(n356) );
  INV_X1 U464 ( .A(n543), .ZN(n372) );
  AND2_X1 U465 ( .A1(n612), .A2(n391), .ZN(n412) );
  NAND2_X1 U466 ( .A1(n628), .A2(n593), .ZN(n368) );
  NAND2_X1 U467 ( .A1(n602), .A2(G469), .ZN(n369) );
  NAND2_X1 U468 ( .A1(n362), .A2(n359), .ZN(n523) );
  XNOR2_X1 U469 ( .A(n360), .B(KEYINPUT87), .ZN(n359) );
  NAND2_X1 U470 ( .A1(n521), .A2(n361), .ZN(n360) );
  NAND2_X1 U471 ( .A1(n609), .A2(KEYINPUT44), .ZN(n361) );
  NAND2_X1 U472 ( .A1(n365), .A2(n364), .ZN(n363) );
  INV_X1 U473 ( .A(n506), .ZN(n364) );
  NAND2_X1 U474 ( .A1(n366), .A2(n354), .ZN(n365) );
  INV_X1 U475 ( .A(n502), .ZN(n366) );
  NAND2_X1 U476 ( .A1(n540), .A2(n678), .ZN(n367) );
  XNOR2_X2 U477 ( .A(n551), .B(n440), .ZN(n665) );
  AND2_X2 U478 ( .A1(n373), .A2(n372), .ZN(n443) );
  NAND2_X1 U479 ( .A1(n373), .A2(n554), .ZN(n673) );
  XNOR2_X2 U480 ( .A(n441), .B(n374), .ZN(n373) );
  NOR2_X2 U481 ( .A1(n579), .A2(n578), .ZN(n581) );
  NOR2_X2 U482 ( .A1(n708), .A2(n599), .ZN(n656) );
  XNOR2_X1 U483 ( .A(KEYINPUT22), .B(n496), .ZN(n500) );
  NOR2_X2 U484 ( .A1(n509), .A2(n497), .ZN(n643) );
  NAND2_X1 U485 ( .A1(n542), .A2(n678), .ZN(n378) );
  XNOR2_X2 U486 ( .A(G143), .B(G128), .ZN(n485) );
  XNOR2_X2 U487 ( .A(n387), .B(G122), .ZN(n475) );
  NOR2_X1 U488 ( .A1(n389), .A2(n661), .ZN(n495) );
  NOR2_X1 U489 ( .A1(n673), .A2(n389), .ZN(n511) );
  XNOR2_X2 U490 ( .A(n465), .B(n464), .ZN(n389) );
  OR2_X1 U491 ( .A1(n692), .A2(n466), .ZN(n393) );
  OR2_X2 U492 ( .A1(n515), .A2(n466), .ZN(n395) );
  NAND2_X1 U493 ( .A1(n692), .A2(n397), .ZN(n396) );
  AND2_X1 U494 ( .A1(n350), .A2(n466), .ZN(n397) );
  XNOR2_X2 U495 ( .A(n443), .B(n442), .ZN(n692) );
  XNOR2_X1 U496 ( .A(n523), .B(n522), .ZN(n597) );
  INV_X1 U497 ( .A(n446), .ZN(n447) );
  OR2_X1 U498 ( .A1(n700), .A2(G902), .ZN(n398) );
  XOR2_X1 U499 ( .A(KEYINPUT104), .B(n534), .Z(n399) );
  XOR2_X1 U500 ( .A(n694), .B(KEYINPUT118), .Z(n400) );
  XNOR2_X1 U501 ( .A(KEYINPUT73), .B(KEYINPUT48), .ZN(n580) );
  INV_X1 U502 ( .A(KEYINPUT33), .ZN(n442) );
  INV_X1 U503 ( .A(KEYINPUT19), .ZN(n458) );
  INV_X1 U504 ( .A(KEYINPUT83), .ZN(n657) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(n457) );
  BUF_X1 U506 ( .A(n597), .Z(n708) );
  XNOR2_X1 U507 ( .A(n412), .B(n411), .ZN(n512) );
  INV_X1 U508 ( .A(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U509 ( .A(n402), .B(KEYINPUT72), .ZN(n403) );
  XNOR2_X1 U510 ( .A(n404), .B(G113), .ZN(n444) );
  XOR2_X1 U511 ( .A(G137), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U512 ( .A(G119), .B(G116), .ZN(n405) );
  XNOR2_X1 U513 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U514 ( .A(n444), .B(n407), .Z(n409) );
  NOR2_X1 U515 ( .A1(G953), .A2(G237), .ZN(n469) );
  NAND2_X1 U516 ( .A1(n469), .A2(G210), .ZN(n408) );
  XNOR2_X1 U517 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U518 ( .A(n439), .B(n410), .ZN(n612) );
  XNOR2_X1 U519 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n413) );
  XNOR2_X1 U520 ( .A(G140), .B(G137), .ZN(n432) );
  XNOR2_X1 U521 ( .A(n474), .B(n432), .ZN(n721) );
  XNOR2_X1 U522 ( .A(n414), .B(KEYINPUT85), .ZN(n418) );
  NAND2_X1 U523 ( .A1(G234), .A2(n526), .ZN(n416) );
  NAND2_X1 U524 ( .A1(n490), .A2(G221), .ZN(n422) );
  XOR2_X1 U525 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n420) );
  XOR2_X2 U526 ( .A(G119), .B(G110), .Z(n446) );
  XNOR2_X1 U527 ( .A(G128), .B(n446), .ZN(n419) );
  XNOR2_X1 U528 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U529 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U530 ( .A(n721), .B(n423), .ZN(n704) );
  NOR2_X1 U531 ( .A1(n704), .A2(G902), .ZN(n427) );
  NAND2_X1 U532 ( .A1(n593), .A2(G234), .ZN(n424) );
  XNOR2_X1 U533 ( .A(n424), .B(KEYINPUT20), .ZN(n428) );
  NAND2_X1 U534 ( .A1(n428), .A2(G217), .ZN(n425) );
  NAND2_X1 U535 ( .A1(n428), .A2(G221), .ZN(n429) );
  XNOR2_X1 U536 ( .A(n429), .B(KEYINPUT21), .ZN(n661) );
  INV_X1 U537 ( .A(n661), .ZN(n430) );
  NAND2_X1 U538 ( .A1(n526), .A2(G227), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n431), .B(KEYINPUT78), .ZN(n433) );
  XNOR2_X1 U540 ( .A(n433), .B(n432), .ZN(n437) );
  XNOR2_X1 U541 ( .A(G110), .B(G107), .ZN(n434) );
  XNOR2_X1 U542 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U543 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U544 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n440) );
  NAND2_X1 U545 ( .A1(n666), .A2(n665), .ZN(n441) );
  OR2_X1 U546 ( .A1(G237), .A2(G902), .ZN(n454) );
  NAND2_X1 U547 ( .A1(G214), .A2(n454), .ZN(n678) );
  XOR2_X1 U548 ( .A(G116), .B(G107), .Z(n486) );
  XNOR2_X1 U549 ( .A(n444), .B(n486), .ZN(n450) );
  NAND2_X1 U550 ( .A1(G224), .A2(n526), .ZN(n451) );
  NAND2_X1 U551 ( .A1(n454), .A2(G210), .ZN(n456) );
  NAND2_X1 U552 ( .A1(G234), .A2(G237), .ZN(n459) );
  XNOR2_X1 U553 ( .A(n459), .B(KEYINPUT14), .ZN(n460) );
  NAND2_X1 U554 ( .A1(G952), .A2(n460), .ZN(n691) );
  NOR2_X1 U555 ( .A1(G953), .A2(n691), .ZN(n530) );
  NAND2_X1 U556 ( .A1(G902), .A2(n460), .ZN(n525) );
  XNOR2_X1 U557 ( .A(G898), .B(KEYINPUT89), .ZN(n711) );
  NAND2_X1 U558 ( .A1(G953), .A2(n711), .ZN(n714) );
  NOR2_X1 U559 ( .A1(n525), .A2(n714), .ZN(n461) );
  NOR2_X1 U560 ( .A1(n530), .A2(n461), .ZN(n462) );
  XNOR2_X1 U561 ( .A(n462), .B(KEYINPUT90), .ZN(n463) );
  NOR2_X2 U562 ( .A1(n535), .A2(n463), .ZN(n465) );
  INV_X1 U563 ( .A(KEYINPUT0), .ZN(n464) );
  XNOR2_X1 U564 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n480) );
  XOR2_X1 U565 ( .A(KEYINPUT11), .B(KEYINPUT94), .Z(n468) );
  XNOR2_X1 U566 ( .A(G131), .B(KEYINPUT93), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n473) );
  XOR2_X1 U568 ( .A(G140), .B(KEYINPUT12), .Z(n471) );
  NAND2_X1 U569 ( .A1(G214), .A2(n469), .ZN(n470) );
  XNOR2_X1 U570 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n473), .B(n472), .ZN(n479) );
  INV_X1 U572 ( .A(n474), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n475), .B(n476), .ZN(n478) );
  XNOR2_X1 U574 ( .A(n481), .B(G475), .ZN(n517) );
  XOR2_X1 U575 ( .A(KEYINPUT9), .B(KEYINPUT96), .Z(n483) );
  XNOR2_X1 U576 ( .A(n483), .B(n482), .ZN(n489) );
  XOR2_X1 U577 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n484) );
  XOR2_X1 U578 ( .A(n485), .B(n484), .Z(n487) );
  XNOR2_X1 U579 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U580 ( .A(n489), .B(n488), .Z(n492) );
  NAND2_X1 U581 ( .A1(G217), .A2(n490), .ZN(n491) );
  XNOR2_X1 U582 ( .A(n492), .B(n491), .ZN(n700) );
  XNOR2_X1 U583 ( .A(G478), .B(n398), .ZN(n516) );
  INV_X1 U584 ( .A(n516), .ZN(n494) );
  NOR2_X1 U585 ( .A1(n609), .A2(KEYINPUT44), .ZN(n502) );
  AND2_X1 U586 ( .A1(n494), .A2(n517), .ZN(n681) );
  NAND2_X1 U587 ( .A1(n681), .A2(n495), .ZN(n496) );
  OR2_X1 U588 ( .A1(n500), .A2(n665), .ZN(n509) );
  INV_X1 U589 ( .A(n531), .ZN(n662) );
  NAND2_X1 U590 ( .A1(n512), .A2(n662), .ZN(n497) );
  XNOR2_X1 U591 ( .A(n665), .B(KEYINPUT88), .ZN(n545) );
  NAND2_X1 U592 ( .A1(n498), .A2(n543), .ZN(n499) );
  NOR2_X1 U593 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U594 ( .A(n501), .B(KEYINPUT32), .ZN(n737) );
  INV_X1 U595 ( .A(KEYINPUT65), .ZN(n507) );
  INV_X1 U596 ( .A(KEYINPUT44), .ZN(n503) );
  NOR2_X1 U597 ( .A1(n503), .A2(KEYINPUT65), .ZN(n504) );
  NAND2_X1 U598 ( .A1(n543), .A2(n531), .ZN(n508) );
  NOR2_X1 U599 ( .A1(n509), .A2(n508), .ZN(n633) );
  XNOR2_X1 U600 ( .A(KEYINPUT31), .B(KEYINPUT92), .ZN(n510) );
  XNOR2_X1 U601 ( .A(n511), .B(n510), .ZN(n652) );
  NAND2_X1 U602 ( .A1(n666), .A2(n551), .ZN(n513) );
  NOR2_X1 U603 ( .A1(n554), .A2(n513), .ZN(n514) );
  NAND2_X1 U604 ( .A1(n350), .A2(n514), .ZN(n637) );
  NAND2_X1 U605 ( .A1(n652), .A2(n637), .ZN(n519) );
  NAND2_X1 U606 ( .A1(n517), .A2(n516), .ZN(n651) );
  XOR2_X1 U607 ( .A(KEYINPUT98), .B(n651), .Z(n588) );
  INV_X1 U608 ( .A(n588), .ZN(n518) );
  OR2_X1 U609 ( .A1(n517), .A2(n516), .ZN(n541) );
  NAND2_X1 U610 ( .A1(n518), .A2(n541), .ZN(n683) );
  AND2_X1 U611 ( .A1(n519), .A2(n683), .ZN(n520) );
  NOR2_X1 U612 ( .A1(n633), .A2(n520), .ZN(n521) );
  NOR2_X2 U613 ( .A1(n597), .A2(n593), .ZN(n524) );
  XNOR2_X1 U614 ( .A(n524), .B(KEYINPUT86), .ZN(n592) );
  XNOR2_X1 U615 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n539) );
  INV_X1 U616 ( .A(n683), .ZN(n538) );
  OR2_X1 U617 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U618 ( .A(KEYINPUT101), .B(n527), .Z(n528) );
  NOR2_X1 U619 ( .A1(G900), .A2(n528), .ZN(n529) );
  NOR2_X1 U620 ( .A1(n530), .A2(n529), .ZN(n556) );
  OR2_X1 U621 ( .A1(n531), .A2(n661), .ZN(n532) );
  NOR2_X1 U622 ( .A1(n556), .A2(n532), .ZN(n542) );
  AND2_X1 U623 ( .A1(n542), .A2(n554), .ZN(n533) );
  XNOR2_X1 U624 ( .A(n533), .B(KEYINPUT28), .ZN(n534) );
  INV_X1 U625 ( .A(n535), .ZN(n536) );
  NAND2_X1 U626 ( .A1(n536), .A2(n551), .ZN(n537) );
  OR2_X1 U627 ( .A1(n399), .A2(n537), .ZN(n647) );
  NOR2_X1 U628 ( .A1(n538), .A2(n647), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n539), .A2(n570), .ZN(n569) );
  INV_X1 U630 ( .A(n574), .ZN(n586) );
  NOR2_X1 U631 ( .A1(n586), .A2(n582), .ZN(n544) );
  XNOR2_X1 U632 ( .A(KEYINPUT36), .B(n544), .ZN(n546) );
  NAND2_X1 U633 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U634 ( .A(n547), .B(KEYINPUT107), .ZN(n732) );
  NAND2_X1 U635 ( .A1(n677), .A2(n678), .ZN(n549) );
  XOR2_X1 U636 ( .A(KEYINPUT106), .B(n549), .Z(n682) );
  NAND2_X1 U637 ( .A1(n682), .A2(n681), .ZN(n550) );
  XNOR2_X1 U638 ( .A(n550), .B(KEYINPUT41), .ZN(n693) );
  INV_X1 U639 ( .A(n551), .ZN(n558) );
  NOR2_X1 U640 ( .A1(n399), .A2(n558), .ZN(n552) );
  NAND2_X1 U641 ( .A1(n693), .A2(n552), .ZN(n553) );
  XOR2_X1 U642 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n565) );
  NAND2_X1 U643 ( .A1(n678), .A2(n554), .ZN(n555) );
  XNOR2_X1 U644 ( .A(KEYINPUT30), .B(n555), .ZN(n562) );
  INV_X1 U645 ( .A(n556), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n666), .A2(n557), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n560), .B(KEYINPUT77), .ZN(n561) );
  NOR2_X1 U648 ( .A1(n562), .A2(n561), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n572), .A2(n677), .ZN(n563) );
  XNOR2_X2 U650 ( .A(n563), .B(KEYINPUT39), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n589), .A2(n634), .ZN(n564) );
  NAND2_X1 U652 ( .A1(n735), .A2(n734), .ZN(n566) );
  XNOR2_X1 U653 ( .A(n566), .B(KEYINPUT46), .ZN(n567) );
  NAND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n579) );
  INV_X1 U655 ( .A(n570), .ZN(n571) );
  NAND2_X1 U656 ( .A1(KEYINPUT47), .A2(n571), .ZN(n576) );
  AND2_X1 U657 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n572), .A2(n575), .ZN(n646) );
  NAND2_X1 U659 ( .A1(n576), .A2(n646), .ZN(n577) );
  XNOR2_X1 U660 ( .A(KEYINPUT84), .B(n577), .ZN(n578) );
  XNOR2_X1 U661 ( .A(n581), .B(n580), .ZN(n591) );
  XNOR2_X1 U662 ( .A(KEYINPUT102), .B(n582), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n583), .A2(n665), .ZN(n585) );
  XNOR2_X1 U664 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n584) );
  XNOR2_X1 U665 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n655) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n654) );
  NAND2_X1 U668 ( .A1(n655), .A2(n654), .ZN(n590) );
  NOR2_X2 U669 ( .A1(n591), .A2(n590), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n592), .A2(n722), .ZN(n596) );
  INV_X1 U671 ( .A(n593), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(KEYINPUT2), .ZN(n595) );
  INV_X1 U673 ( .A(n598), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n656), .A2(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U675 ( .A1(n703), .A2(G469), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n601) );
  XNOR2_X1 U677 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U678 ( .A(G952), .ZN(n605) );
  NOR2_X2 U679 ( .A1(n606), .A2(n707), .ZN(n608) );
  INV_X1 U680 ( .A(KEYINPUT119), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n608), .B(n607), .ZN(G54) );
  XOR2_X1 U682 ( .A(n351), .B(G122), .Z(G24) );
  NAND2_X1 U683 ( .A1(n703), .A2(G472), .ZN(n614) );
  XNOR2_X1 U684 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(KEYINPUT62), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X2 U687 ( .A1(n615), .A2(n707), .ZN(n617) );
  INV_X1 U688 ( .A(KEYINPUT63), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(G57) );
  NAND2_X1 U690 ( .A1(n703), .A2(G475), .ZN(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT67), .B(KEYINPUT120), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT59), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U694 ( .A1(n623), .A2(n707), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n624) );
  XOR2_X1 U696 ( .A(n624), .B(KEYINPUT68), .Z(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(G60) );
  NAND2_X1 U698 ( .A1(n703), .A2(G210), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n352), .B(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U702 ( .A1(n631), .A2(n707), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U704 ( .A(G101), .B(n633), .Z(G3) );
  NOR2_X1 U705 ( .A1(n541), .A2(n637), .ZN(n635) );
  XOR2_X1 U706 ( .A(G104), .B(n635), .Z(n636) );
  XNOR2_X1 U707 ( .A(KEYINPUT110), .B(n636), .ZN(G6) );
  NOR2_X1 U708 ( .A1(n651), .A2(n637), .ZN(n642) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n639) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT111), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U712 ( .A(KEYINPUT26), .B(n640), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G9) );
  XOR2_X1 U714 ( .A(G110), .B(n643), .Z(G12) );
  NOR2_X1 U715 ( .A1(n651), .A2(n647), .ZN(n645) );
  XNOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G30) );
  XNOR2_X1 U718 ( .A(G143), .B(n646), .ZN(G45) );
  NOR2_X1 U719 ( .A1(n541), .A2(n647), .ZN(n648) );
  XOR2_X1 U720 ( .A(G146), .B(n648), .Z(G48) );
  NOR2_X1 U721 ( .A1(n652), .A2(n541), .ZN(n650) );
  XNOR2_X1 U722 ( .A(G113), .B(KEYINPUT113), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(G15) );
  NOR2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U725 ( .A(G116), .B(n653), .Z(G18) );
  XNOR2_X1 U726 ( .A(G134), .B(n654), .ZN(G36) );
  XNOR2_X1 U727 ( .A(G140), .B(n655), .ZN(G42) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n697) );
  XOR2_X1 U730 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n664) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n672) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U736 ( .A(KEYINPUT115), .B(n669), .Z(n670) );
  NOR2_X1 U737 ( .A1(n670), .A2(n554), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NAND2_X1 U741 ( .A1(n693), .A2(n676), .ZN(n688) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(KEYINPUT117), .B(n679), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n692), .A2(n686), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U749 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  NOR2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U754 ( .A1(n703), .A2(G478), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n707), .A2(n702), .ZN(G63) );
  NAND2_X1 U757 ( .A1(n703), .A2(G217), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n707), .A2(n706), .ZN(G66) );
  NOR2_X1 U760 ( .A1(n708), .A2(G953), .ZN(n713) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n709) );
  XOR2_X1 U762 ( .A(KEYINPUT61), .B(n709), .Z(n710) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n719) );
  XOR2_X1 U765 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n717) );
  NAND2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n720), .B(n721), .ZN(n726) );
  XNOR2_X1 U770 ( .A(n722), .B(n726), .ZN(n723) );
  XNOR2_X1 U771 ( .A(KEYINPUT124), .B(n723), .ZN(n724) );
  NOR2_X1 U772 ( .A1(G953), .A2(n724), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n725), .B(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U774 ( .A(n726), .B(G227), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G900), .ZN(n728) );
  XNOR2_X1 U776 ( .A(KEYINPUT126), .B(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G125), .B(n732), .ZN(n733) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U781 ( .A(n734), .B(G131), .ZN(G33) );
  XOR2_X1 U782 ( .A(G137), .B(n735), .Z(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT127), .B(n736), .ZN(G39) );
  XOR2_X1 U784 ( .A(n737), .B(G119), .Z(G21) );
endmodule

