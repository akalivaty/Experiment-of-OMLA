//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT94), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G15gat), .ZN(new_n208));
  INV_X1    g007(.A(G15gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G22gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n210), .A3(new_n205), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n203), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n210), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(new_n205), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n202), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n202), .A3(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G29gat), .A2(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT15), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT15), .A4(new_n226), .ZN(new_n230));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n230), .A2(new_n231), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n232), .B2(new_n234), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n219), .B(new_n220), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n234), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n212), .A2(new_n202), .A3(new_n217), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n218), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n242), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247));
  INV_X1    g046(.A(new_n240), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n220), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n239), .B(KEYINPUT13), .Z(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  AOI211_X1 g052(.A(KEYINPUT95), .B(new_n253), .C1(new_n249), .C2(new_n242), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n245), .B(new_n246), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT93), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n266), .B(KEYINPUT86), .Z(new_n267));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269));
  INV_X1    g068(.A(G141gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G148gat), .ZN(new_n271));
  INV_X1    g070(.A(G148gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G141gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n273), .A3(KEYINPUT79), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n270), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n276), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT80), .B(G155gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT2), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n275), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  INV_X1    g083(.A(G211gat), .ZN(new_n285));
  INV_X1    g084(.A(G218gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n284), .C1(KEYINPUT22), .C2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(KEYINPUT87), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(KEYINPUT22), .B2(new_n287), .ZN(new_n291));
  INV_X1    g090(.A(new_n283), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n289), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n282), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G155gat), .B(G162gat), .Z(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(KEYINPUT2), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n277), .A3(new_n268), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n269), .B1(new_n279), .B2(G162gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n297), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n294), .B1(new_n304), .B2(new_n290), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n267), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n293), .B2(new_n288), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n308), .A2(KEYINPUT88), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n297), .B1(new_n308), .B2(KEYINPUT88), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n305), .A2(new_n266), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n207), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G78gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n313), .A3(new_n207), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  OAI21_X1  g118(.A(G78gat), .B1(new_n319), .B2(new_n314), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT31), .B(G50gat), .ZN(new_n321));
  INV_X1    g120(.A(G106gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n318), .B2(new_n320), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT35), .ZN(new_n328));
  INV_X1    g127(.A(new_n294), .ZN(new_n329));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n335));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n339), .B1(new_n349), .B2(KEYINPUT66), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(G183gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT67), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n347), .A2(G190gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n332), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n344), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n346), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n344), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n370));
  AND2_X1   g169(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n342), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n340), .A2(new_n341), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(KEYINPUT65), .C1(new_n371), .C2(new_n370), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n368), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n331), .B1(new_n379), .B2(new_n290), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n330), .B1(new_n368), .B2(new_n378), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n329), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n368), .B2(new_n378), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n383), .B(new_n294), .C1(new_n331), .C2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n390), .B2(KEYINPUT78), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n389), .B1(new_n382), .B2(new_n385), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n327), .A2(new_n328), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT32), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n377), .A2(KEYINPUT25), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT67), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT67), .B1(new_n352), .B2(new_n353), .ZN(new_n400));
  INV_X1    g199(.A(new_n360), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT66), .B1(new_n349), .B2(new_n357), .ZN(new_n403));
  AOI21_X1  g202(.A(G190gat), .B1(new_n352), .B2(new_n351), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT28), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n367), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n346), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n409));
  INV_X1    g208(.A(G113gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G120gat), .ZN(new_n411));
  INV_X1    g210(.A(G120gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G113gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G134gat), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT1), .B1(new_n416), .B2(G127gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n418));
  INV_X1    g217(.A(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G134gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G127gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n425), .A3(G134gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n419), .B2(G134gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n416), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT70), .A4(G134gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT1), .B1(new_n411), .B2(new_n413), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n409), .B(new_n422), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n430), .A3(new_n431), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT69), .B(G127gat), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT70), .B1(new_n440), .B2(G134gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n422), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT72), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI22_X1  g243(.A1(new_n398), .A2(new_n408), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n443), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n409), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(KEYINPUT72), .A3(new_n443), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n368), .A4(new_n378), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G227gat), .ZN(new_n451));
  INV_X1    g250(.A(G233gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n397), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G15gat), .B(G43gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT73), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT33), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT74), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n445), .B2(new_n449), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n463));
  INV_X1    g262(.A(new_n459), .ZN(new_n464));
  NOR4_X1   g263(.A1(new_n462), .A2(new_n463), .A3(new_n397), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n462), .A2(KEYINPUT33), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n458), .B1(new_n462), .B2(new_n397), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n460), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n449), .A3(new_n461), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(KEYINPUT75), .A2(KEYINPUT34), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  OAI221_X1 g274(.A(new_n473), .B1(new_n466), .B2(new_n467), .C1(new_n460), .C2(new_n465), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n423), .A2(new_n425), .A3(G134gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n432), .B1(new_n479), .B2(KEYINPUT70), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n436), .B1(new_n480), .B2(new_n428), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n307), .B1(new_n481), .B2(new_n422), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n282), .A2(new_n443), .A3(new_n442), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n478), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n447), .A2(KEYINPUT4), .A3(new_n282), .A4(new_n448), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n446), .A2(new_n492), .A3(new_n304), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n493), .A3(new_n485), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n487), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n447), .A2(new_n282), .A3(new_n448), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n490), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n493), .A2(new_n478), .A3(new_n485), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n485), .A3(new_n493), .A4(new_n491), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n499), .B1(new_n496), .B2(new_n490), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n505), .A2(new_n487), .B1(new_n506), .B2(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT91), .ZN(new_n508));
  XNOR2_X1  g307(.A(G57gat), .B(G85gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT82), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G1gat), .B(G29gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n504), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n507), .B2(new_n514), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n514), .B1(new_n495), .B2(new_n501), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n516), .A2(new_n519), .B1(new_n520), .B2(new_n518), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n396), .A2(new_n477), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n501), .A3(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n517), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT84), .B1(new_n526), .B2(new_n520), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n515), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n517), .A4(new_n525), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n520), .A2(new_n518), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n524), .B1(new_n532), .B2(new_n395), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n326), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n324), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n477), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n524), .A3(new_n395), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n515), .B1(new_n507), .B2(KEYINPUT91), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n502), .A2(new_n503), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n519), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n382), .A2(new_n385), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT37), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  INV_X1    g346(.A(new_n389), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n382), .A2(new_n385), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n544), .A2(new_n531), .A3(new_n390), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n551), .A2(new_n390), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n521), .A2(new_n555), .A3(KEYINPUT92), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT38), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT39), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  AOI211_X1 g360(.A(new_n561), .B(new_n485), .C1(new_n506), .C2(new_n493), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n497), .A2(new_n500), .A3(new_n493), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT89), .B1(new_n563), .B2(new_n486), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n446), .A2(new_n492), .A3(new_n304), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n499), .B(new_n566), .C1(new_n496), .C2(new_n490), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n561), .B1(new_n567), .B2(new_n485), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(KEYINPUT89), .A3(new_n486), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n484), .A2(new_n486), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(new_n560), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n565), .A2(new_n572), .A3(new_n514), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT40), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(KEYINPUT90), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n516), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n395), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n559), .A2(new_n327), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT36), .B1(new_n477), .B2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584));
  AOI211_X1 g383(.A(new_n583), .B(new_n584), .C1(new_n475), .C2(new_n476), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n532), .A2(new_n524), .A3(new_n395), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n536), .B1(new_n587), .B2(new_n533), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n581), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n265), .B1(new_n541), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n237), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n594), .A2(KEYINPUT8), .ZN(new_n595));
  NOR2_X1   g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(KEYINPUT8), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT98), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n601), .A2(new_n603), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n600), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT98), .B1(new_n598), .B2(new_n599), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n602), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n592), .A2(new_n235), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n611), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n248), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n591), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n236), .B2(new_n237), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n603), .B1(new_n601), .B2(new_n610), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n602), .B(new_n609), .C1(new_n597), .C2(new_n600), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n240), .ZN(new_n626));
  INV_X1    g425(.A(new_n591), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n622), .A2(new_n626), .A3(new_n618), .A4(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n620), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT99), .A3(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(G57gat), .A2(G64gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G71gat), .A2(G78gat), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT9), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G57gat), .A2(G64gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n644));
  INV_X1    g443(.A(new_n639), .ZN(new_n645));
  NOR2_X1   g444(.A1(G71gat), .A2(G78gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G71gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n316), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(KEYINPUT96), .A3(new_n639), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  INV_X1    g451(.A(new_n642), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n637), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n652), .A2(new_n654), .A3(KEYINPUT96), .A4(new_n641), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT21), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n219), .A2(new_n220), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n219), .A2(new_n220), .A3(new_n657), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G231gat), .A2(G233gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n656), .B2(KEYINPUT21), .ZN(new_n666));
  XNOR2_X1  g465(.A(G127gat), .B(G155gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT97), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT21), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n655), .A3(new_n670), .A4(new_n664), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n669), .B1(new_n666), .B2(new_n671), .ZN(new_n674));
  XOR2_X1   g473(.A(G183gat), .B(G211gat), .Z(new_n675));
  NOR3_X1   g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n666), .A2(new_n671), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n668), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n663), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n675), .B1(new_n673), .B2(new_n674), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n677), .A3(new_n672), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n662), .A4(new_n660), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n633), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n621), .A2(new_n628), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n621), .A2(new_n628), .A3(KEYINPUT100), .A4(new_n686), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n636), .A2(new_n685), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(new_n656), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n623), .B2(new_n624), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n615), .A2(new_n611), .A3(new_n656), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G230gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n452), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT10), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n697), .A2(new_n698), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n656), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n695), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(G120gat), .B(G148gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(G176gat), .B(G204gat), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n709), .B(new_n710), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n695), .B(new_n711), .C1(new_n703), .C2(new_n707), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n694), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n590), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n532), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(G1gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1324gat));
  XNOR2_X1  g520(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n722));
  INV_X1    g521(.A(new_n395), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n590), .A2(new_n723), .A3(new_n717), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT16), .B(G8gat), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT105), .Z(new_n726));
  OAI21_X1  g525(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(G8gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n727), .B(new_n728), .C1(new_n724), .C2(new_n730), .ZN(G1325gat));
  OAI21_X1  g530(.A(new_n209), .B1(new_n718), .B2(new_n477), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n586), .A2(new_n209), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n718), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g535(.A1(new_n718), .A2(new_n327), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT43), .B(G22gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1327gat));
  AND2_X1   g538(.A1(new_n689), .A2(new_n690), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n636), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n685), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n590), .A2(new_n715), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n532), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n221), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n559), .A2(new_n327), .A3(new_n580), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n588), .A2(new_n586), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT109), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n581), .A2(new_n753), .A3(new_n586), .A4(new_n588), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n749), .B1(new_n755), .B2(new_n541), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n541), .A2(new_n589), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n748), .B1(new_n757), .B2(new_n741), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n715), .B(KEYINPUT108), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n265), .A3(new_n685), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G29gat), .B1(new_n763), .B2(new_n532), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n764), .ZN(G1328gat));
  NAND3_X1  g564(.A1(new_n744), .A2(new_n222), .A3(new_n723), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT46), .Z(new_n767));
  OAI21_X1  g566(.A(G36gat), .B1(new_n763), .B2(new_n395), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1329gat));
  INV_X1    g568(.A(new_n586), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n770), .B(new_n762), .C1(new_n756), .C2(new_n758), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G43gat), .ZN(new_n772));
  INV_X1    g571(.A(G43gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n477), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n744), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1330gat));
  OAI211_X1 g579(.A(new_n536), .B(new_n762), .C1(new_n756), .C2(new_n758), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G50gat), .ZN(new_n782));
  INV_X1    g581(.A(G50gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n744), .A2(new_n783), .A3(new_n536), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n786), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(new_n788), .A3(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1331gat));
  AND2_X1   g589(.A1(new_n588), .A2(new_n586), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n753), .B1(new_n791), .B2(new_n581), .ZN(new_n792));
  INV_X1    g591(.A(new_n754), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n541), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n255), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n261), .B1(new_n255), .B2(KEYINPUT93), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n694), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n794), .A2(new_n795), .A3(new_n761), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n522), .B1(KEYINPUT35), .B2(new_n539), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n752), .B2(new_n754), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n761), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT111), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n745), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g606(.A(KEYINPUT49), .B(G64gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n723), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n800), .A2(new_n804), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n810), .A2(new_n395), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1333gat));
  NAND3_X1  g611(.A1(new_n800), .A2(new_n770), .A3(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G71gat), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n800), .A2(new_n648), .A3(new_n804), .A4(new_n774), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(KEYINPUT50), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1334gat));
  NOR2_X1   g619(.A1(new_n810), .A2(new_n327), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(new_n316), .ZN(G1335gat));
  NOR3_X1   g621(.A1(new_n798), .A2(new_n715), .A3(new_n685), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n759), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G85gat), .B1(new_n824), .B2(new_n532), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n743), .A2(new_n265), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n794), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n802), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(new_n605), .A3(new_n745), .A4(new_n716), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n825), .A2(new_n832), .ZN(G1336gat));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n723), .B(new_n823), .C1(new_n756), .C2(new_n758), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G92gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n395), .A2(G92gat), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n761), .B(new_n838), .C1(new_n828), .C2(new_n830), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AND4_X1   g640(.A1(new_n835), .A2(new_n837), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n836), .B2(G92gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n835), .B1(new_n843), .B2(new_n839), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(G1337gat));
  XNOR2_X1  g644(.A(KEYINPUT113), .B(G99gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n774), .A3(new_n716), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n586), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n846), .ZN(G1338gat));
  OAI211_X1 g648(.A(new_n536), .B(new_n823), .C1(new_n756), .C2(new_n758), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G106gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n327), .A2(G106gat), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n761), .B(new_n852), .C1(new_n828), .C2(new_n830), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1339gat));
  NAND3_X1  g657(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n705), .A2(new_n706), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n702), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n705), .A2(KEYINPUT115), .A3(new_n706), .A4(new_n701), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT54), .A4(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n711), .B1(new_n707), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(KEYINPUT55), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n863), .B(new_n711), .C1(new_n699), .C2(new_n702), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT55), .B1(new_n865), .B2(new_n867), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n250), .A2(new_n251), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n239), .B1(new_n238), .B2(new_n242), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n260), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n255), .A2(new_n262), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n872), .A2(new_n741), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n255), .B2(new_n262), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n715), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n872), .B2(new_n798), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n880), .B2(new_n741), .ZN(new_n881));
  INV_X1    g680(.A(new_n685), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n693), .A2(new_n883), .A3(new_n265), .A4(new_n715), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n740), .A2(new_n692), .A3(new_n685), .A4(new_n636), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n265), .A3(new_n886), .A4(new_n715), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT114), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n881), .A2(new_n882), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n532), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n537), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n395), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n410), .B1(new_n892), .B2(new_n265), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n889), .A2(new_n536), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n745), .A2(new_n395), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n477), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(G113gat), .A3(new_n798), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT116), .Z(G1340gat));
  NAND3_X1  g699(.A1(new_n891), .A2(new_n395), .A3(new_n716), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n760), .A2(new_n412), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n901), .A2(new_n412), .B1(new_n897), .B2(new_n902), .ZN(G1341gat));
  INV_X1    g702(.A(new_n897), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n882), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n685), .A2(new_n440), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n905), .A2(new_n440), .B1(new_n892), .B2(new_n906), .ZN(G1342gat));
  OAI21_X1  g706(.A(G134gat), .B1(new_n904), .B2(new_n742), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n723), .A2(G134gat), .A3(new_n742), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n908), .A2(new_n909), .B1(new_n891), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n909), .A3(new_n910), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n891), .A2(KEYINPUT117), .A3(new_n909), .A4(new_n910), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n911), .B2(new_n916), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1343gat));
  NOR2_X1   g719(.A1(new_n770), .A2(new_n327), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n890), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n395), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n270), .B1(new_n924), .B2(new_n265), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n889), .B2(new_n327), .ZN(new_n927));
  INV_X1    g726(.A(new_n871), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n869), .A3(new_n868), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n265), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n742), .B1(new_n930), .B2(new_n879), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n685), .B1(new_n931), .B2(new_n877), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n887), .B(new_n883), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT57), .B(new_n536), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n770), .A2(new_n895), .ZN(new_n937));
  INV_X1    g736(.A(new_n889), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n938), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n536), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n265), .A2(new_n270), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n925), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n936), .A2(new_n716), .A3(new_n937), .A4(new_n939), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n272), .A2(KEYINPUT59), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n881), .A2(new_n882), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n887), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT57), .B1(new_n953), .B2(new_n536), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n938), .A2(new_n956), .A3(KEYINPUT57), .A4(new_n536), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n937), .A2(new_n716), .ZN(new_n959));
  OAI21_X1  g758(.A(G148gat), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n949), .A2(new_n951), .B1(KEYINPUT59), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n923), .A2(new_n272), .A3(new_n395), .A4(new_n716), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n945), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(KEYINPUT59), .ZN(new_n965));
  INV_X1    g764(.A(new_n951), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n950), .B1(new_n946), .B2(new_n947), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(KEYINPUT122), .A3(new_n962), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n964), .A2(new_n969), .ZN(G1345gat));
  OAI21_X1  g769(.A(new_n279), .B1(new_n940), .B2(new_n882), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n882), .A2(new_n279), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n924), .B2(new_n972), .ZN(G1346gat));
  OAI21_X1  g772(.A(G162gat), .B1(new_n940), .B2(new_n742), .ZN(new_n974));
  OR4_X1    g773(.A1(G162gat), .A2(new_n922), .A3(new_n723), .A4(new_n742), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1347gat));
  NAND2_X1  g775(.A1(new_n723), .A2(new_n532), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(new_n477), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n894), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(G169gat), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(new_n265), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n889), .A2(new_n745), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n536), .A2(new_n395), .A3(new_n477), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n798), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n981), .B1(new_n980), .B2(new_n986), .ZN(G1348gat));
  AOI21_X1  g786(.A(G176gat), .B1(new_n985), .B2(new_n716), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n894), .A2(G176gat), .A3(new_n761), .A4(new_n978), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(G1349gat));
  OAI21_X1  g791(.A(G183gat), .B1(new_n979), .B2(new_n882), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n685), .A2(new_n358), .A3(new_n359), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n984), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g795(.A1(new_n985), .A2(new_n339), .A3(new_n741), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  OAI21_X1  g797(.A(G190gat), .B1(new_n979), .B2(new_n742), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT61), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1351gat));
  INV_X1    g800(.A(new_n958), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n770), .A2(new_n977), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(G197gat), .B1(new_n1004), .B2(new_n265), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n770), .A2(new_n395), .A3(new_n327), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n982), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n1007), .A2(G197gat), .A3(new_n265), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1005), .A2(new_n1009), .ZN(G1352gat));
  NOR3_X1   g809(.A1(new_n1007), .A2(G204gat), .A3(new_n715), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT62), .ZN(new_n1012));
  OAI21_X1  g811(.A(KEYINPUT126), .B1(new_n1004), .B2(new_n760), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G204gat), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n1004), .A2(KEYINPUT126), .A3(new_n760), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1353gat));
  OAI21_X1  g815(.A(G211gat), .B1(new_n1004), .B2(new_n882), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n1017), .A2(KEYINPUT63), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(KEYINPUT63), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1007), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1020), .A2(new_n285), .A3(new_n685), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1022), .ZN(G1354gat));
  OAI21_X1  g822(.A(G218gat), .B1(new_n1004), .B2(new_n742), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1020), .A2(new_n286), .A3(new_n741), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1024), .A2(new_n1025), .ZN(G1355gat));
endmodule


