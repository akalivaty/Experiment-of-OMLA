//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n463), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n472), .A2(new_n473), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n498), .B(new_n499), .C1(new_n473), .C2(new_n472), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n466), .B2(new_n498), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n494), .B(new_n496), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n506), .B(KEYINPUT5), .C1(new_n507), .C2(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(KEYINPUT71), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT71), .B1(new_n511), .B2(G543), .ZN(new_n512));
  OAI211_X1 g087(.A(G62), .B(new_n508), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n505), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(G651), .ZN(new_n523));
  AND4_X1   g098(.A1(G50), .A2(new_n522), .A3(G543), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n513), .B2(new_n514), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(KEYINPUT75), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT73), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n520), .A2(new_n521), .B1(new_n519), .B2(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT5), .B1(new_n506), .B2(new_n507), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n506), .B1(new_n507), .B2(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n530), .A2(new_n531), .A3(new_n534), .A4(new_n508), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT74), .B(G88), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n517), .A2(new_n526), .A3(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  AND2_X1   g114(.A1(new_n529), .A2(new_n535), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT76), .B(G89), .Z(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(G76), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n516), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n530), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G51), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G63), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n528), .A2(new_n549), .B1(new_n543), .B2(new_n544), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n548), .B1(G651), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n542), .A2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  NAND2_X1  g128(.A1(new_n540), .A2(G90), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n534), .A2(G64), .A3(new_n508), .ZN(new_n555));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n516), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(KEYINPUT77), .B1(G52), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  NAND2_X1  g137(.A1(new_n540), .A2(G81), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n528), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n558), .B2(G43), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n529), .A2(new_n535), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT78), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n529), .A2(new_n578), .A3(G91), .A4(new_n535), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT79), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n528), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(KEYINPUT80), .A3(G651), .ZN(new_n588));
  INV_X1    g163(.A(G53), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT9), .B1(new_n546), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n558), .A2(new_n591), .A3(G53), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n587), .A2(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n580), .A2(new_n593), .ZN(G299));
  INV_X1    g169(.A(G74), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n516), .B1(new_n528), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(G49), .B2(new_n558), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n529), .A2(G87), .A3(new_n535), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n528), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n558), .B2(G48), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n529), .A2(G86), .A3(new_n535), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n540), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n528), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(G47), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n609), .A2(G651), .B1(new_n558), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n606), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n575), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT82), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n528), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(new_n558), .B2(G54), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT83), .Z(G148));
  NOR2_X1   g208(.A1(new_n569), .A2(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n624), .A2(new_n631), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n466), .A2(new_n464), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n488), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n490), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n463), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n643), .A2(new_n644), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT86), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2451), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n657), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2454), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n642), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n650), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT91), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n697), .B(new_n696), .S(new_n689), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n704), .B(new_n705), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n702), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n686), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(new_n709), .A3(new_n685), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(KEYINPUT36), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n717));
  OR2_X1    g292(.A1(G6), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(G305), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT32), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1981), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT94), .B(G16), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G166), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G22), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1971), .ZN(new_n728));
  MUX2_X1   g303(.A(G23), .B(G288), .S(G16), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT33), .B(G1976), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n722), .A2(new_n723), .A3(new_n728), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT92), .B(G29), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n488), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n490), .A2(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n463), .A2(G107), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(new_n743), .B2(new_n733), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT35), .B(G1991), .Z(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  MUX2_X1   g321(.A(G24), .B(G290), .S(new_n725), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1986), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n732), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n727), .B(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n731), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n723), .B1(new_n754), .B2(new_n722), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n717), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n722), .A2(new_n728), .A3(new_n731), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT34), .ZN(new_n758));
  INV_X1    g333(.A(new_n717), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n732), .A4(new_n749), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT99), .B(G28), .Z(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT30), .B2(new_n763), .ZN(new_n765));
  INV_X1    g340(.A(new_n733), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n762), .B(new_n765), .C1(new_n649), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n733), .A2(G27), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n733), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT102), .B(G2078), .Z(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G26), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n733), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n488), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n490), .A2(G128), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G29), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n771), .B1(new_n769), .B2(new_n770), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2090), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n733), .A2(G35), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n492), .B2(new_n766), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT29), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n786), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT103), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n792), .B2(new_n787), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n790), .A2(KEYINPUT103), .A3(G2090), .A4(new_n791), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n724), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n569), .B2(new_n724), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1341), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G21), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G168), .B2(G16), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G1966), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(G1966), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n801), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n719), .A2(G5), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G301), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(G1961), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n798), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G139), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n467), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n463), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n781), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n781), .A2(G33), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT97), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(new_n822), .C1(new_n820), .C2(new_n781), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2072), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n781), .A2(G32), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n488), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n490), .A2(G129), .ZN(new_n831));
  NAND3_X1  g406(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT26), .Z(new_n833));
  AND3_X1   g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n834), .B2(new_n781), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT27), .B(G1996), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(G160), .A2(G29), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT24), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(G34), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(G34), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n766), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G2084), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT98), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n850), .A3(new_n838), .A4(new_n828), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n724), .A2(G20), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT23), .Z(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G299), .B2(G16), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1956), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n812), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n837), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n809), .A2(new_n810), .B1(new_n835), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n845), .B2(new_n846), .ZN(new_n861));
  AOI211_X1 g436(.A(KEYINPUT100), .B(G2084), .C1(new_n840), .C2(new_n844), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(new_n859), .C1(new_n861), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n719), .A2(G4), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n624), .B2(new_n719), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT96), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(new_n867), .C1(new_n624), .C2(new_n719), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(G1348), .ZN(new_n873));
  INV_X1    g448(.A(G1348), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n869), .B2(new_n871), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n864), .B(new_n866), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n857), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n761), .A2(new_n877), .ZN(G311));
  AND3_X1   g453(.A1(new_n761), .A2(KEYINPUT104), .A3(new_n877), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT104), .B1(new_n761), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(G150));
  NAND2_X1  g456(.A1(new_n540), .A2(G93), .ZN(new_n882));
  NAND2_X1  g457(.A1(G80), .A2(G543), .ZN(new_n883));
  INV_X1    g458(.A(G67), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n528), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n885), .A2(G651), .B1(new_n558), .B2(G55), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G860), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n618), .A2(new_n623), .ZN(new_n890));
  OR3_X1    g465(.A1(new_n890), .A2(KEYINPUT105), .A3(new_n631), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT105), .B1(new_n890), .B2(new_n631), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT38), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n563), .A2(new_n882), .A3(new_n567), .A4(new_n886), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n563), .A2(new_n567), .B1(new_n882), .B2(new_n886), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n899), .A3(new_n892), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n894), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n894), .B2(new_n900), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT39), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G860), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n889), .B1(new_n907), .B2(new_n908), .ZN(G145));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(new_n820), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n494), .A2(new_n496), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT107), .B1(new_n501), .B2(new_n502), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n498), .B1(new_n472), .B2(new_n473), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT4), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n500), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n780), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n834), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n834), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n919), .A2(new_n834), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n820), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n488), .A2(G142), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n490), .A2(G130), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n463), .A2(G118), .ZN(new_n929));
  OAI21_X1  g504(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(new_n640), .Z(new_n932));
  XNOR2_X1  g507(.A(new_n743), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n910), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g510(.A(KEYINPUT108), .B(new_n933), .C1(new_n923), .C2(new_n925), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n923), .A2(new_n925), .A3(new_n933), .ZN(new_n938));
  OR2_X1    g513(.A1(G160), .A2(new_n649), .ZN(new_n939));
  NAND2_X1  g514(.A1(G160), .A2(new_n649), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(G162), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  AOI21_X1  g518(.A(G162), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n492), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT110), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT111), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n941), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n923), .A2(new_n925), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n933), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n955), .C1(new_n935), .C2(new_n936), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n958), .B(new_n959), .C1(new_n935), .C2(new_n936), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n942), .A2(new_n944), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n957), .A2(KEYINPUT40), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT40), .B1(new_n957), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(G395));
  NAND2_X1  g540(.A1(new_n624), .A2(new_n628), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n890), .A2(G299), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT41), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n635), .B(new_n898), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n968), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT113), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  XNOR2_X1  g552(.A(G166), .B(G290), .ZN(new_n978));
  XOR2_X1   g553(.A(G288), .B(G305), .Z(new_n979));
  OR2_X1    g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT42), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n976), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n974), .A2(new_n975), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n986), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  OAI21_X1  g563(.A(G868), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G868), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n887), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(G295));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n991), .ZN(G331));
  NAND2_X1  g568(.A1(new_n980), .A2(new_n982), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n568), .A2(new_n887), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n995), .A2(G286), .A3(new_n895), .ZN(new_n996));
  AOI21_X1  g571(.A(G286), .B1(new_n995), .B2(new_n895), .ZN(new_n997));
  OAI21_X1  g572(.A(G301), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G168), .B1(new_n896), .B2(new_n897), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(G286), .A3(new_n895), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(G171), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n968), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n969), .A2(new_n971), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n994), .B(new_n1004), .C1(new_n1005), .C2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(G37), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n969), .A2(new_n1009), .A3(new_n971), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n998), .A2(new_n1001), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n968), .A2(KEYINPUT114), .A3(KEYINPUT41), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n994), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1008), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n968), .B1(new_n998), .B2(new_n1001), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n972), .B2(new_n1011), .ZN(new_n1018));
  AOI21_X1  g593(.A(G37), .B1(new_n1018), .B2(new_n994), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1004), .B1(new_n1005), .B2(new_n1002), .ZN(new_n1020));
  INV_X1    g595(.A(new_n994), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1008), .A2(new_n1014), .A3(KEYINPUT43), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1015), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(G397));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n918), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n494), .A2(new_n496), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n915), .A2(new_n916), .A3(new_n500), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n916), .B1(new_n915), .B2(new_n500), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(KEYINPUT116), .A3(new_n1032), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n915), .A2(new_n500), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT45), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n488), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n477), .B1(new_n476), .B2(G2105), .ZN(new_n1045));
  AOI211_X1 g620(.A(KEYINPUT67), .B(new_n463), .C1(new_n474), .C2(new_n475), .ZN(new_n1046));
  OAI211_X1 g621(.A(G40), .B(new_n1044), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT56), .B(G2072), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1040), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1956), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1047), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1384), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n580), .A2(new_n593), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1050), .A2(KEYINPUT122), .A3(new_n1058), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1061), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1038), .A2(new_n479), .A3(G40), .A4(new_n1056), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G2067), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1053), .B1(new_n503), .B2(new_n1056), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1047), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1038), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1348), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n624), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1067), .A2(new_n1075), .B1(new_n1065), .B2(new_n1059), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n890), .A2(new_n1073), .A3(new_n1069), .A4(KEYINPUT60), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n874), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n890), .C1(G2067), .C2(new_n1068), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1074), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1081), .B2(KEYINPUT60), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1062), .A2(new_n1050), .A3(new_n1064), .A4(new_n1058), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1058), .A2(new_n1050), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT61), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1086), .C1(new_n1067), .C2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n568), .A2(KEYINPUT124), .ZN(new_n1089));
  INV_X1    g664(.A(G1996), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1040), .A2(new_n1090), .A3(new_n1048), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1068), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1091), .A2(KEYINPUT123), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT123), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT59), .B(new_n1089), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1076), .B1(new_n1088), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G8), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n918), .A2(G1384), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1052), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n597), .A2(new_n598), .A3(G1976), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1976), .B1(new_n597), .B2(new_n598), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1104), .B(new_n1107), .C1(KEYINPUT52), .C2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1068), .A2(new_n1106), .A3(G8), .A4(new_n1105), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1068), .A2(G8), .A3(new_n1108), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G305), .A2(G1981), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n603), .B2(new_n604), .ZN(new_n1118));
  OR3_X1    g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1104), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G303), .A2(G8), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1971), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1078), .A2(G2090), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1127), .B(G8), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n479), .B(G40), .C1(new_n1042), .C2(KEYINPUT45), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1134), .A2(G1971), .B1(new_n1078), .B2(G2090), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(KEYINPUT117), .A3(G8), .A4(new_n1127), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1122), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n918), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT116), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1048), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n751), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n787), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1102), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT120), .B1(new_n1144), .B2(new_n1127), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1127), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1140), .A2(new_n751), .B1(new_n1142), .B2(new_n787), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1146), .B(new_n1147), .C1(new_n1148), .C2(new_n1102), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1078), .A2(new_n810), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(G2078), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1044), .A2(G40), .A3(new_n1153), .ZN(new_n1154));
  OAI221_X1 g729(.A(new_n1154), .B1(new_n463), .B2(new_n470), .C1(new_n1103), .C2(KEYINPUT45), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1040), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G2078), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n1134), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(G171), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1140), .B2(G2078), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT45), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n503), .A2(new_n1032), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n479), .A2(new_n1163), .A3(G40), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(new_n1153), .B1(new_n1078), .B2(new_n810), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(G301), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1160), .A2(KEYINPUT54), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(G1966), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1071), .A2(new_n1072), .A3(new_n846), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(G168), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(G8), .ZN(new_n1173));
  AOI21_X1  g748(.A(G168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT51), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT51), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(new_n1176), .A3(G8), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AND4_X1   g753(.A1(new_n1137), .A2(new_n1150), .A3(new_n1168), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1157), .A2(new_n1159), .A3(G171), .ZN(new_n1181));
  AOI21_X1  g756(.A(G301), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT125), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1185), .B(new_n1180), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1101), .A2(new_n1179), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G286), .A2(new_n1102), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1150), .A2(new_n1137), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1189), .A2(KEYINPUT63), .A3(new_n1190), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1135), .A2(G8), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1147), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1137), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1194), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(G288), .A2(G1976), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT119), .Z(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1120), .B2(new_n1119), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1104), .B1(new_n1205), .B2(new_n1115), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1206), .B1(new_n1207), .B2(new_n1122), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1175), .A2(new_n1209), .A3(new_n1177), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1182), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1150), .A2(new_n1137), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1188), .A2(new_n1202), .A3(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1103), .A2(KEYINPUT45), .A3(new_n1047), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n742), .B(new_n745), .ZN(new_n1218));
  NAND2_X1  g793(.A1(G290), .A2(G1986), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n834), .B(G1996), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n780), .B(G2067), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1218), .A2(new_n1219), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(G290), .A2(G1986), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1225), .B(KEYINPUT115), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1217), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1216), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1226), .A2(KEYINPUT48), .A3(new_n1217), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1217), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(KEYINPUT48), .B1(new_n1226), .B2(new_n1217), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1221), .A2(new_n834), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n1217), .ZN(new_n1236));
  XOR2_X1   g811(.A(new_n1236), .B(KEYINPUT126), .Z(new_n1237));
  NAND2_X1  g812(.A1(new_n1217), .A2(new_n1090), .ZN(new_n1238));
  XOR2_X1   g813(.A(new_n1238), .B(KEYINPUT46), .Z(new_n1239));
  NOR2_X1   g814(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1240), .B(KEYINPUT47), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n780), .A2(new_n783), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n743), .A2(new_n745), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1242), .B1(new_n1243), .B2(new_n1222), .ZN(new_n1244));
  AOI211_X1 g819(.A(new_n1234), .B(new_n1241), .C1(new_n1217), .C2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1228), .A2(new_n1245), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g821(.A1(G227), .A2(new_n461), .ZN(new_n1248));
  XOR2_X1   g822(.A(new_n1248), .B(KEYINPUT127), .Z(new_n1249));
  NOR2_X1   g823(.A1(G401), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g824(.A1(new_n712), .A2(new_n714), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1251), .B1(new_n957), .B2(new_n962), .ZN(new_n1252));
  AND2_X1   g826(.A1(new_n1013), .A2(new_n1004), .ZN(new_n1253));
  OAI211_X1 g827(.A(new_n1019), .B(new_n1015), .C1(new_n1253), .C2(new_n994), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1018), .A2(new_n994), .ZN(new_n1255));
  OAI21_X1  g829(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g830(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  AND2_X1   g831(.A1(new_n1252), .A2(new_n1257), .ZN(G308));
  NAND2_X1  g832(.A1(new_n1252), .A2(new_n1257), .ZN(G225));
endmodule


