//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n463), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n468), .A2(new_n469), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n466), .A2(new_n470), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n491), .B(KEYINPUT71), .C1(new_n469), .C2(new_n468), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT71), .B1(new_n476), .B2(new_n491), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n484), .B2(G126), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n511), .A2(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n509), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n515), .A2(new_n516), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n529), .A2(G51), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  INV_X1    g111(.A(G77), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n522), .A2(new_n536), .B1(new_n537), .B2(new_n528), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n540), .B1(new_n537), .B2(new_n528), .C1(new_n522), .C2(new_n536), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(G651), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT75), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n539), .A2(new_n544), .A3(new_n541), .A4(G651), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n511), .A2(new_n546), .B1(new_n517), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n543), .A2(new_n545), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT77), .B(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n511), .A2(new_n553), .B1(new_n517), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n555), .B1(KEYINPUT76), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n562), .B(G651), .C1(new_n557), .C2(new_n559), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n552), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n517), .ZN(new_n565));
  INV_X1    g140(.A(new_n554), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n529), .B2(G43), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n559), .B1(new_n506), .B2(G56), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT76), .B1(new_n568), .B2(new_n508), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n567), .A2(new_n569), .A3(new_n563), .A4(new_n552), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT80), .Z(G188));
  NAND2_X1  g154(.A1(new_n517), .A2(KEYINPUT81), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n506), .A2(new_n510), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(G91), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n529), .B2(G53), .ZN(new_n585));
  INV_X1    g160(.A(G53), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g163(.A1(new_n514), .A2(new_n513), .A3(KEYINPUT82), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n504), .B2(new_n505), .ZN(new_n591));
  OAI21_X1  g166(.A(G65), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G78), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n508), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G299));
  OR2_X1    g171(.A1(new_n506), .A2(G74), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n529), .B2(G49), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n580), .A2(G87), .A3(new_n582), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n522), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n529), .B2(G48), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n580), .A2(G86), .A3(new_n582), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(G85), .A2(new_n565), .B1(new_n529), .B2(G47), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n508), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n580), .A2(G92), .A3(new_n582), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n580), .A2(KEYINPUT10), .A3(G92), .A4(new_n582), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n529), .A2(G54), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G66), .B1(new_n589), .B2(new_n591), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G651), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n615), .A2(KEYINPUT83), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT83), .B1(new_n615), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n595), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n630), .B2(G860), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT84), .Z(G148));
  NAND2_X1  g207(.A1(new_n615), .A2(new_n621), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n615), .A2(new_n621), .A3(KEYINPUT83), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n572), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g215(.A1(new_n466), .A2(new_n470), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n474), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT12), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n644), .A3(new_n474), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n482), .A2(G135), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n484), .A2(G123), .ZN(new_n652));
  OR2_X1    g227(.A1(G99), .A2(G2105), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n653), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n647), .B2(new_n648), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(new_n657), .ZN(G156));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  INV_X1    g237(.A(G2435), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT15), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G2435), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G2438), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(G2438), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n662), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n674));
  INV_X1    g249(.A(new_n662), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(G2438), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT14), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n669), .A2(new_n671), .A3(new_n662), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n661), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n673), .B2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n660), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1341), .B(G1348), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n684), .A2(new_n660), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n682), .B(new_n661), .C1(new_n673), .C2(new_n680), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2451), .B(G2454), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n689), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G14), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n689), .B2(new_n693), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n659), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n689), .A2(new_n693), .ZN(new_n700));
  INV_X1    g275(.A(new_n695), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n702), .A2(KEYINPUT89), .A3(G14), .A4(new_n696), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G401));
  INV_X1    g280(.A(KEYINPUT18), .ZN(new_n706));
  XOR2_X1   g281(.A(G2084), .B(G2090), .Z(new_n707));
  XNOR2_X1  g282(.A(G2067), .B(G2678), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT17), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT90), .B(G2100), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(G2072), .B(G2078), .Z(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n709), .B2(KEYINPUT18), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G2096), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n714), .B(new_n717), .ZN(G227));
  XOR2_X1   g293(.A(G1991), .B(G1996), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1971), .B(G1976), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT19), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(G1956), .B(G2474), .Z(new_n724));
  XOR2_X1   g299(.A(G1961), .B(G1966), .Z(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n723), .A2(new_n726), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT20), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n732), .B(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n738), .B2(new_n730), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n720), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(G1981), .B(G1986), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n735), .A2(new_n739), .A3(new_n720), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n742), .ZN(new_n745));
  INV_X1    g320(.A(new_n743), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n740), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(G229));
  XOR2_X1   g324(.A(KEYINPUT33), .B(G1976), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G23), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(G288), .B2(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(G6), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G305), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT32), .B(G1981), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n751), .A2(new_n755), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n751), .B2(new_n755), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n754), .A2(G22), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G166), .B2(new_n754), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G1971), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n757), .A2(new_n759), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n763), .A2(G1971), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT34), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n482), .A2(G131), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G119), .ZN(new_n774));
  OR2_X1    g349(.A1(G95), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n772), .B1(new_n778), .B2(new_n771), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT35), .B(G1991), .Z(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  MUX2_X1   g356(.A(G24), .B(G290), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n781), .B(new_n783), .C1(KEYINPUT93), .C2(KEYINPUT36), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n769), .A2(new_n770), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n785), .B(new_n786), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n482), .A2(G141), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n484), .A2(G129), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n474), .A2(G105), .ZN(new_n790));
  NAND3_X1  g365(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT26), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n771), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n771), .B2(G32), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT97), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n771), .A2(G27), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT101), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n771), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n799), .B1(G2078), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n754), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n754), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G1966), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n771), .A2(G26), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(G128), .A2(new_n484), .B1(new_n482), .B2(G140), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT95), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n810), .B1(new_n817), .B2(new_n771), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G2067), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n805), .A2(G1966), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT30), .B(G28), .ZN(new_n821));
  OR2_X1    g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  NAND2_X1  g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(new_n771), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n655), .B2(new_n771), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n807), .A2(new_n819), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n771), .A2(G33), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n466), .A2(new_n470), .A3(G127), .ZN(new_n828));
  NAND2_X1  g403(.A1(G115), .A2(G2104), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n463), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G139), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n477), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n827), .B1(new_n836), .B2(new_n771), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(G2072), .Z(new_n838));
  XOR2_X1   g413(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n754), .A2(G20), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n595), .B2(new_n754), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1956), .Z(new_n843));
  NAND4_X1  g418(.A1(new_n803), .A2(new_n826), .A3(new_n838), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n771), .A2(G35), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G162), .B2(new_n771), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT29), .Z(new_n847));
  INV_X1    g422(.A(G2090), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n802), .A2(G2078), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT24), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n771), .B1(new_n852), .B2(G34), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(G34), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G160), .B2(G29), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(G2084), .ZN(new_n856));
  NOR4_X1   g431(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n572), .A2(new_n754), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n754), .B2(G19), .ZN(new_n859));
  INV_X1    g434(.A(G1341), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NOR2_X1   g437(.A1(G5), .A2(G16), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT99), .Z(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(G301), .B2(new_n754), .ZN(new_n865));
  INV_X1    g440(.A(G1961), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n857), .A2(new_n861), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n796), .A2(new_n797), .B1(G2084), .B2(new_n855), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n866), .B2(new_n865), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT100), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n844), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n754), .A2(G4), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n624), .B2(new_n754), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT94), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G1348), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n787), .A2(new_n872), .A3(new_n876), .ZN(G150));
  INV_X1    g452(.A(G150), .ZN(G311));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(G860), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n508), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT103), .B(G55), .ZN(new_n883));
  INV_X1    g458(.A(G93), .ZN(new_n884));
  OAI22_X1  g459(.A1(new_n511), .A2(new_n883), .B1(new_n517), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n564), .B2(new_n571), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n567), .A2(new_n563), .A3(new_n569), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT38), .ZN(new_n893));
  INV_X1    g468(.A(new_n624), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n630), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(KEYINPUT78), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n886), .B1(new_n896), .B2(new_n570), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(new_n890), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(G559), .A3(new_n624), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n880), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT104), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n906), .A3(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n902), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n887), .A2(G860), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n879), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n907), .A2(new_n905), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT106), .B(new_n911), .C1(new_n914), .C2(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G145));
  NAND2_X1  g491(.A1(new_n794), .A2(new_n836), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n793), .B1(new_n830), .B2(new_n835), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n482), .A2(G142), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n484), .A2(G130), .ZN(new_n921));
  OR2_X1    g496(.A1(G106), .A2(G2105), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n922), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n643), .A2(new_n645), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n643), .B2(new_n645), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n925), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n918), .B(new_n917), .C1(new_n929), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n816), .A2(new_n502), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n816), .A2(new_n502), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n778), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n817), .A2(G164), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n777), .A3(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(G160), .A2(new_n655), .ZN(new_n940));
  NAND2_X1  g515(.A1(G160), .A2(new_n655), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(G162), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n928), .A2(new_n930), .A3(new_n935), .A4(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n939), .B2(new_n944), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT40), .Z(G395));
  INV_X1    g525(.A(G288), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(G303), .ZN(new_n952));
  XNOR2_X1  g527(.A(G290), .B(G305), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G299), .A2(new_n633), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n595), .B1(new_n615), .B2(new_n621), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n637), .A2(KEYINPUT107), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n635), .A2(new_n965), .A3(new_n630), .A4(new_n636), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n964), .A2(new_n898), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n898), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n624), .B2(new_n630), .ZN(new_n970));
  INV_X1    g545(.A(new_n966), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n892), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n898), .A3(new_n966), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT41), .B1(new_n961), .B2(new_n962), .ZN(new_n974));
  INV_X1    g549(.A(new_n633), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n595), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT41), .ZN(new_n977));
  NAND2_X1  g552(.A1(G299), .A2(new_n633), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(KEYINPUT108), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n963), .C1(new_n967), .C2(new_n968), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n960), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n960), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(G868), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n886), .A2(G868), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(G295));
  INV_X1    g565(.A(G868), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n984), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n959), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n960), .A2(new_n982), .A3(new_n984), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n995), .B2(new_n988), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n997), .A3(new_n989), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(G331));
  NAND3_X1  g574(.A1(new_n963), .A2(KEYINPUT112), .A3(new_n977), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n979), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1002), .A3(new_n974), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n526), .A2(new_n533), .A3(KEYINPUT111), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n532), .A2(new_n531), .ZN(new_n1006));
  INV_X1    g581(.A(G51), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n511), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1008), .B2(new_n525), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n548), .B1(new_n542), .B2(KEYINPUT75), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n545), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n545), .B2(new_n1011), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1013), .A2(new_n1014), .B1(new_n897), .B2(new_n890), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G301), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n888), .A2(new_n1017), .A3(new_n891), .A4(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1003), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n963), .A3(new_n1018), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n954), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n979), .A2(new_n974), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1015), .A2(new_n963), .A3(new_n1018), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n954), .ZN(new_n1027));
  AOI21_X1  g602(.A(G37), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT43), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n954), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(KEYINPUT44), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n1029), .B2(KEYINPUT43), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1027), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1019), .A2(new_n980), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1027), .A3(new_n1021), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n946), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1036), .A2(new_n1039), .A3(KEYINPUT43), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1031), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1034), .A2(new_n1035), .B1(KEYINPUT44), .B2(new_n1042), .ZN(G397));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n604), .A2(new_n1044), .A3(new_n605), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G48), .ZN(new_n1047));
  INV_X1    g622(.A(G86), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n511), .A2(new_n1047), .B1(new_n517), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  OAI221_X1 g626(.A(new_n1051), .B1(new_n517), .B2(new_n1048), .C1(new_n1047), .C2(new_n511), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n603), .A2(G651), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(G1981), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1049), .A2(KEYINPUT114), .B1(G651), .B2(new_n603), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1044), .B1(new_n1057), .B2(new_n1052), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1045), .A2(KEYINPUT115), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  INV_X1    g637(.A(G40), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n473), .A2(new_n1063), .A3(new_n479), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1384), .B1(new_n497), .B2(new_n501), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1056), .B(new_n1067), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1061), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G288), .A2(G1976), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1046), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(new_n1066), .B(KEYINPUT116), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n951), .A2(G1976), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n951), .A2(G1976), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1074), .A2(KEYINPUT52), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1069), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n479), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n471), .A2(new_n472), .ZN(new_n1080));
  OAI211_X1 g655(.A(G40), .B(new_n1079), .C1(new_n1080), .C2(new_n463), .ZN(new_n1081));
  INV_X1    g656(.A(G1384), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n502), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1083), .B2(KEYINPUT50), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1065), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n848), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1971), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1065), .A2(KEYINPUT45), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1064), .B1(new_n1065), .B2(KEYINPUT45), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1062), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT55), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1071), .A2(new_n1072), .B1(new_n1078), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1069), .A2(new_n1077), .A3(new_n1076), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(KEYINPUT118), .C1(new_n1096), .C2(new_n1093), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1078), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G2084), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1084), .A2(new_n1104), .A3(new_n1086), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1062), .B(G286), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1097), .A2(new_n1108), .A3(KEYINPUT63), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT45), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1081), .B1(new_n1083), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1971), .B1(new_n1112), .B2(new_n1089), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1064), .B1(new_n1065), .B2(new_n1085), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1086), .A2(KEYINPUT117), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1065), .A2(new_n1116), .A3(new_n1085), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n848), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1095), .B1(new_n1119), .B2(new_n1062), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1099), .A2(new_n1120), .A3(new_n1097), .A4(new_n1108), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1098), .B1(new_n1110), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1105), .A2(new_n1107), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G168), .A2(new_n1062), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1129), .A3(G168), .ZN(new_n1133));
  AND2_X1   g708(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1126), .A2(G8), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1125), .B(new_n1132), .C1(new_n1135), .C2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1133), .A2(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT62), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1099), .A2(new_n1097), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1120), .ZN(new_n1144));
  INV_X1    g719(.A(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1112), .A2(new_n1145), .A3(new_n1089), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n866), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1112), .A2(KEYINPUT53), .A3(new_n1145), .A4(new_n1089), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(G171), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1143), .A2(new_n1144), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1139), .A2(new_n1142), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1083), .B2(new_n1081), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1064), .A2(new_n1065), .A3(KEYINPUT120), .ZN(new_n1159));
  AOI21_X1  g734(.A(G2067), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1348), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n633), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT56), .B(G2072), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1112), .A2(new_n1089), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1118), .B2(G1956), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n595), .B(KEYINPUT57), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1163), .A2(new_n1164), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT121), .B1(new_n1162), .B2(new_n633), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1168), .B(new_n1166), .C1(new_n1118), .C2(G1956), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1170), .A2(new_n1171), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1160), .ZN(new_n1178));
  INV_X1    g753(.A(G1348), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1150), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1183), .A3(new_n975), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n633), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT58), .B(G1341), .Z(new_n1188));
  NAND3_X1  g763(.A1(new_n1158), .A2(new_n1159), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(G1996), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1112), .A2(new_n1190), .A3(new_n1089), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1187), .B1(new_n1192), .B2(new_n572), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1192), .A2(new_n572), .A3(new_n1187), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1184), .B(new_n1185), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1196), .A2(KEYINPUT61), .A3(new_n1172), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1176), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1196), .B1(new_n1199), .B2(new_n1174), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1177), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1090), .A2(new_n1091), .A3(G2078), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1204), .A2(KEYINPUT53), .B1(new_n1150), .B2(new_n866), .ZN(new_n1205));
  AOI21_X1  g780(.A(G301), .B1(new_n1205), .B2(new_n1148), .ZN(new_n1206));
  AND4_X1   g781(.A1(G301), .A2(new_n1148), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT54), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1205), .A2(G301), .A3(new_n1148), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT54), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1154), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1212), .B(new_n1213), .C1(new_n1141), .C2(new_n1140), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n1124), .B(new_n1156), .C1(new_n1203), .C2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1081), .A2(new_n1065), .A3(KEYINPUT45), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n816), .A2(G2067), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n816), .A2(G2067), .ZN(new_n1218));
  AND2_X1   g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n793), .B(new_n1190), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n778), .A2(new_n780), .ZN(new_n1221));
  OR2_X1    g796(.A1(new_n778), .A2(new_n780), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(G290), .B(G1986), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1216), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1215), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1216), .A2(new_n1190), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT46), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1219), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1216), .B1(new_n1229), .B2(new_n793), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1231), .B(KEYINPUT47), .Z(new_n1232));
  NAND2_X1  g807(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1217), .B1(new_n1233), .B2(new_n1221), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1216), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT125), .Z(new_n1236));
  NOR2_X1   g811(.A1(G290), .A2(G1986), .ZN(new_n1237));
  AOI21_X1  g812(.A(KEYINPUT48), .B1(new_n1216), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g813(.A1(new_n1216), .A2(KEYINPUT48), .A3(new_n1237), .ZN(new_n1239));
  AOI211_X1 g814(.A(new_n1238), .B(new_n1239), .C1(new_n1216), .C2(new_n1223), .ZN(new_n1240));
  NOR3_X1   g815(.A1(new_n1232), .A2(new_n1236), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1226), .A2(new_n1241), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g817(.A(new_n748), .B1(new_n947), .B2(new_n948), .ZN(new_n1244));
  NOR2_X1   g818(.A1(G227), .A2(new_n461), .ZN(new_n1245));
  INV_X1    g819(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g820(.A(new_n1246), .B1(new_n699), .B2(new_n703), .ZN(new_n1247));
  AOI21_X1  g821(.A(new_n1244), .B1(new_n1247), .B2(KEYINPUT126), .ZN(new_n1248));
  NAND2_X1  g822(.A1(new_n704), .A2(new_n1245), .ZN(new_n1249));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g824(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1253));
  NOR3_X1   g827(.A1(new_n1042), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1247), .A2(KEYINPUT126), .ZN(new_n1255));
  AOI211_X1 g829(.A(new_n1250), .B(new_n1246), .C1(new_n699), .C2(new_n703), .ZN(new_n1256));
  NOR3_X1   g830(.A1(new_n1255), .A2(new_n1256), .A3(new_n1244), .ZN(new_n1257));
  NAND3_X1  g831(.A1(new_n1023), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1258));
  NAND3_X1  g832(.A1(new_n1032), .A2(new_n1038), .A3(new_n946), .ZN(new_n1259));
  NAND2_X1  g833(.A1(new_n1259), .A2(KEYINPUT43), .ZN(new_n1260));
  NAND2_X1  g834(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g835(.A(KEYINPUT127), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g836(.A1(new_n1254), .A2(new_n1262), .ZN(G308));
  OAI21_X1  g837(.A(new_n1253), .B1(new_n1042), .B2(new_n1252), .ZN(new_n1264));
  NAND3_X1  g838(.A1(new_n1257), .A2(new_n1261), .A3(KEYINPUT127), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n1264), .A2(new_n1265), .ZN(G225));
endmodule


