

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605;

  NOR2_X1 U330 ( .A1(n603), .A2(n569), .ZN(n472) );
  XNOR2_X1 U331 ( .A(n394), .B(n393), .ZN(n478) );
  INV_X1 U332 ( .A(n598), .ZN(n569) );
  INV_X1 U333 ( .A(n547), .ZN(n541) );
  INV_X1 U334 ( .A(n525), .ZN(n538) );
  XNOR2_X2 U335 ( .A(G197GAT), .B(G218GAT), .ZN(n368) );
  XNOR2_X2 U336 ( .A(n369), .B(n368), .ZN(n381) );
  BUF_X1 U337 ( .A(n509), .Z(n298) );
  NOR2_X1 U338 ( .A1(n424), .A2(n423), .ZN(n425) );
  XNOR2_X1 U339 ( .A(n363), .B(n362), .ZN(n525) );
  XNOR2_X1 U340 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n367) );
  AND2_X1 U341 ( .A1(n397), .A2(n536), .ZN(n545) );
  XOR2_X1 U342 ( .A(n374), .B(n373), .Z(n299) );
  XOR2_X1 U343 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n300) );
  INV_X1 U344 ( .A(G1GAT), .ZN(n339) );
  XNOR2_X1 U345 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U346 ( .A(n370), .B(n311), .ZN(n312) );
  XNOR2_X1 U347 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U348 ( .A(n441), .B(n312), .ZN(n313) );
  XNOR2_X1 U349 ( .A(n375), .B(n299), .ZN(n376) );
  NOR2_X1 U350 ( .A1(n525), .A2(n481), .ZN(n588) );
  XNOR2_X1 U351 ( .A(n377), .B(n376), .ZN(n379) );
  NOR2_X1 U352 ( .A1(n547), .A2(n485), .ZN(n584) );
  INV_X1 U353 ( .A(G183GAT), .ZN(n487) );
  XOR2_X1 U354 ( .A(n594), .B(KEYINPUT41), .Z(n578) );
  XOR2_X1 U355 ( .A(KEYINPUT105), .B(n463), .Z(n509) );
  XNOR2_X1 U356 ( .A(n487), .B(KEYINPUT124), .ZN(n488) );
  XNOR2_X1 U357 ( .A(n464), .B(G29GAT), .ZN(n465) );
  XNOR2_X1 U358 ( .A(n489), .B(n488), .ZN(G1350GAT) );
  XNOR2_X1 U359 ( .A(n466), .B(n465), .ZN(G1328GAT) );
  NAND2_X1 U360 ( .A1(G230GAT), .A2(G233GAT), .ZN(n306) );
  XOR2_X1 U361 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n302) );
  XNOR2_X1 U362 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n304) );
  XOR2_X1 U364 ( .A(G120GAT), .B(KEYINPUT75), .Z(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U367 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n308) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G92GAT), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(G85GAT), .B(n309), .Z(n441) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n310), .B(G148GAT), .ZN(n370) );
  XOR2_X1 U373 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n311) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n319) );
  XOR2_X1 U375 ( .A(G64GAT), .B(KEYINPUT76), .Z(n316) );
  XNOR2_X1 U376 ( .A(G176GAT), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n388) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G57GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n317), .B(KEYINPUT13), .ZN(n444) );
  XNOR2_X1 U380 ( .A(n388), .B(n444), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n594) );
  XOR2_X1 U382 ( .A(G15GAT), .B(G113GAT), .Z(n321) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G197GAT), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n323) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n337) );
  XOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT69), .Z(n456) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G141GAT), .Z(n327) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U393 ( .A(n456), .B(n328), .Z(n330) );
  NAND2_X1 U394 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U396 ( .A(n331), .B(KEYINPUT70), .Z(n335) );
  XOR2_X1 U397 ( .A(G29GAT), .B(G43GAT), .Z(n333) );
  XNOR2_X1 U398 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n430) );
  XNOR2_X1 U400 ( .A(n430), .B(KEYINPUT30), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n574) );
  INV_X1 U403 ( .A(n574), .ZN(n589) );
  OR2_X1 U404 ( .A1(n594), .A2(n589), .ZN(n493) );
  XNOR2_X1 U405 ( .A(KEYINPUT88), .B(KEYINPUT1), .ZN(n338) );
  XNOR2_X1 U406 ( .A(n300), .B(n338), .ZN(n342) );
  NAND2_X1 U407 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XOR2_X1 U408 ( .A(n343), .B(KEYINPUT92), .Z(n350) );
  XOR2_X1 U409 ( .A(G134GAT), .B(KEYINPUT78), .Z(n427) );
  XOR2_X1 U410 ( .A(n427), .B(G162GAT), .Z(n347) );
  XOR2_X1 U411 ( .A(G120GAT), .B(KEYINPUT80), .Z(n345) );
  XNOR2_X1 U412 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n401) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(n401), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n348), .B(KEYINPUT4), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U418 ( .A(G85GAT), .B(G155GAT), .Z(n352) );
  XNOR2_X1 U419 ( .A(G127GAT), .B(G148GAT), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U421 ( .A(n354), .B(n353), .Z(n363) );
  XOR2_X1 U422 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n356) );
  XNOR2_X1 U423 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U425 ( .A(G141GAT), .B(n357), .ZN(n378) );
  INV_X1 U426 ( .A(n378), .ZN(n361) );
  XOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT89), .Z(n359) );
  XNOR2_X1 U428 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U431 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n365) );
  NAND2_X1 U432 ( .A1(G228GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U434 ( .A(n366), .B(KEYINPUT83), .Z(n372) );
  INV_X1 U435 ( .A(n367), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n381), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U438 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XOR2_X1 U439 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XNOR2_X1 U440 ( .A(n438), .B(n443), .ZN(n375) );
  XOR2_X1 U441 ( .A(G204GAT), .B(G211GAT), .Z(n374) );
  XNOR2_X1 U442 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n482) );
  XOR2_X1 U444 ( .A(n482), .B(KEYINPUT28), .Z(n542) );
  NOR2_X1 U445 ( .A1(n538), .A2(n542), .ZN(n397) );
  INV_X1 U446 ( .A(KEYINPUT94), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n383) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n385) );
  INV_X1 U450 ( .A(KEYINPUT93), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U452 ( .A(G36GAT), .B(G190GAT), .Z(n426) );
  XOR2_X1 U453 ( .A(n426), .B(G92GAT), .Z(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U456 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n391) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n398) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(G183GAT), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n392), .B(G211GAT), .ZN(n448) );
  XNOR2_X1 U461 ( .A(n398), .B(n448), .ZN(n393) );
  INV_X1 U462 ( .A(KEYINPUT95), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n478), .B(n395), .ZN(n396) );
  XNOR2_X1 U464 ( .A(KEYINPUT27), .B(n396), .ZN(n536) );
  XNOR2_X1 U465 ( .A(n545), .B(KEYINPUT96), .ZN(n414) );
  XOR2_X1 U466 ( .A(G15GAT), .B(G127GAT), .Z(n455) );
  XOR2_X1 U467 ( .A(n398), .B(n455), .Z(n400) );
  XNOR2_X1 U468 ( .A(G134GAT), .B(G190GAT), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U470 ( .A(n401), .B(KEYINPUT20), .Z(n403) );
  NAND2_X1 U471 ( .A1(G227GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U473 ( .A(n405), .B(n404), .Z(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT82), .B(KEYINPUT65), .Z(n407) );
  XNOR2_X1 U475 ( .A(G43GAT), .B(G99GAT), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U477 ( .A(G71GAT), .B(G176GAT), .Z(n409) );
  XNOR2_X1 U478 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n547) );
  NAND2_X1 U482 ( .A1(n414), .A2(n547), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n415), .B(KEYINPUT97), .ZN(n424) );
  NAND2_X1 U484 ( .A1(n478), .A2(n541), .ZN(n416) );
  NAND2_X1 U485 ( .A1(n482), .A2(n416), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n417), .B(KEYINPUT25), .ZN(n421) );
  NOR2_X1 U487 ( .A1(n482), .A2(n541), .ZN(n419) );
  XOR2_X1 U488 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n418) );
  XOR2_X1 U489 ( .A(n419), .B(n418), .Z(n587) );
  AND2_X1 U490 ( .A1(n587), .A2(n536), .ZN(n420) );
  NOR2_X1 U491 ( .A1(n421), .A2(n420), .ZN(n422) );
  NOR2_X1 U492 ( .A1(n525), .A2(n422), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n425), .B(KEYINPUT99), .ZN(n491) );
  XOR2_X1 U494 ( .A(KEYINPUT64), .B(n426), .Z(n429) );
  XNOR2_X1 U495 ( .A(G218GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U497 ( .A(G106GAT), .B(n430), .Z(n432) );
  NAND2_X1 U498 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U500 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U501 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n436) );
  XNOR2_X1 U502 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n435) );
  XNOR2_X1 U503 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U504 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n572) );
  XNOR2_X1 U507 ( .A(KEYINPUT36), .B(n572), .ZN(n603) );
  XOR2_X1 U508 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U509 ( .A1(G231GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U511 ( .A(n447), .B(KEYINPUT12), .Z(n450) );
  XNOR2_X1 U512 ( .A(n448), .B(KEYINPUT15), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n452) );
  XNOR2_X1 U515 ( .A(G78GAT), .B(G64GAT), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U517 ( .A(n454), .B(n453), .Z(n458) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n598) );
  NOR2_X1 U520 ( .A1(n603), .A2(n598), .ZN(n459) );
  AND2_X1 U521 ( .A1(n491), .A2(n459), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT37), .ZN(n524) );
  OR2_X1 U523 ( .A1(n493), .A2(n524), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n461) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n298), .A2(n525), .ZN(n466) );
  XOR2_X1 U527 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n464) );
  XNOR2_X1 U528 ( .A(n598), .B(KEYINPUT115), .ZN(n555) );
  XOR2_X1 U529 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n484) );
  XNOR2_X1 U530 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n467), .B(KEYINPUT118), .ZN(n480) );
  INV_X1 U532 ( .A(n572), .ZN(n583) );
  NAND2_X1 U533 ( .A1(n574), .A2(n578), .ZN(n468) );
  XNOR2_X1 U534 ( .A(KEYINPUT46), .B(n468), .ZN(n469) );
  NAND2_X1 U535 ( .A1(n469), .A2(n555), .ZN(n470) );
  NOR2_X1 U536 ( .A1(n583), .A2(n470), .ZN(n471) );
  XNOR2_X1 U537 ( .A(KEYINPUT47), .B(n471), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT45), .B(n472), .Z(n473) );
  NOR2_X1 U539 ( .A1(n594), .A2(n473), .ZN(n474) );
  NAND2_X1 U540 ( .A1(n589), .A2(n474), .ZN(n475) );
  NAND2_X1 U541 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n477), .B(KEYINPUT48), .ZN(n549) );
  BUF_X1 U543 ( .A(n478), .Z(n527) );
  AND2_X1 U544 ( .A1(n549), .A2(n527), .ZN(n479) );
  XNOR2_X1 U545 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U546 ( .A1(n588), .A2(n482), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U548 ( .A(n584), .ZN(n486) );
  NOR2_X1 U549 ( .A1(n555), .A2(n486), .ZN(n489) );
  NOR2_X1 U550 ( .A1(n583), .A2(n569), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT16), .ZN(n492) );
  NAND2_X1 U552 ( .A1(n492), .A2(n491), .ZN(n512) );
  NOR2_X1 U553 ( .A1(n493), .A2(n512), .ZN(n502) );
  NAND2_X1 U554 ( .A1(n502), .A2(n525), .ZN(n497) );
  XOR2_X1 U555 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n495) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U559 ( .A1(n502), .A2(n527), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U562 ( .A1(n502), .A2(n541), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G15GAT), .B(n501), .ZN(G1326GAT) );
  XOR2_X1 U565 ( .A(G22GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U566 ( .A1(n502), .A2(n542), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n298), .A2(n527), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U571 ( .A1(n298), .A2(n541), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U574 ( .A1(n298), .A2(n542), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT108), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  NAND2_X1 U577 ( .A1(n578), .A2(n589), .ZN(n523) );
  NOR2_X1 U578 ( .A1(n523), .A2(n512), .ZN(n513) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(n513), .Z(n519) );
  NAND2_X1 U580 ( .A1(n525), .A2(n519), .ZN(n514) );
  XNOR2_X1 U581 ( .A(KEYINPUT42), .B(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n527), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n516), .B(KEYINPUT110), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n541), .A2(n519), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U589 ( .A1(n519), .A2(n542), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n522), .Z(G1335GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n525), .A2(n532), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  XOR2_X1 U598 ( .A(G99GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U599 ( .A1(n532), .A2(n541), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(G1338GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n534) );
  NAND2_X1 U602 ( .A1(n532), .A2(n542), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U604 ( .A(G106GAT), .B(n535), .Z(G1339GAT) );
  INV_X1 U605 ( .A(n549), .ZN(n540) );
  INV_X1 U606 ( .A(n536), .ZN(n537) );
  OR2_X1 U607 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n562) );
  NAND2_X1 U609 ( .A1(n541), .A2(n562), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n542), .A2(KEYINPUT116), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n545), .A2(KEYINPUT116), .ZN(n546) );
  NOR2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n559), .A2(n574), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT49), .Z(n554) );
  NAND2_X1 U619 ( .A1(n578), .A2(n559), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1341GAT) );
  INV_X1 U621 ( .A(n559), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT50), .B(n557), .Z(n558) );
  XNOR2_X1 U624 ( .A(G127GAT), .B(n558), .ZN(G1342GAT) );
  XOR2_X1 U625 ( .A(G134GAT), .B(KEYINPUT51), .Z(n561) );
  NAND2_X1 U626 ( .A1(n583), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1343GAT) );
  NAND2_X1 U628 ( .A1(n587), .A2(n562), .ZN(n571) );
  NOR2_X1 U629 ( .A1(n589), .A2(n571), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1344GAT) );
  INV_X1 U632 ( .A(n578), .ZN(n565) );
  NOR2_X1 U633 ( .A1(n565), .A2(n571), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(G148GAT), .B(n568), .ZN(G1345GAT) );
  NOR2_X1 U637 ( .A1(n569), .A2(n571), .ZN(n570) );
  XOR2_X1 U638 ( .A(G155GAT), .B(n570), .Z(G1346GAT) );
  NOR2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U640 ( .A(G162GAT), .B(n573), .Z(G1347GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n576) );
  NAND2_X1 U642 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(G169GAT), .B(n577), .ZN(G1348GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n580) );
  NAND2_X1 U646 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U648 ( .A(G176GAT), .B(KEYINPUT56), .Z(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(G1349GAT) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(KEYINPUT58), .ZN(n586) );
  XNOR2_X1 U652 ( .A(G190GAT), .B(n586), .ZN(G1351GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n602) );
  NOR2_X1 U654 ( .A1(n589), .A2(n602), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1352GAT) );
  XOR2_X1 U659 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n596) );
  INV_X1 U660 ( .A(n602), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n599), .A2(n594), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U663 ( .A(G204GAT), .B(n597), .ZN(G1353GAT) );
  XOR2_X1 U664 ( .A(G211GAT), .B(KEYINPUT127), .Z(n601) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U666 ( .A(n601), .B(n600), .ZN(G1354GAT) );
  NOR2_X1 U667 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U668 ( .A(KEYINPUT62), .B(n604), .Z(n605) );
  XNOR2_X1 U669 ( .A(G218GAT), .B(n605), .ZN(G1355GAT) );
endmodule

