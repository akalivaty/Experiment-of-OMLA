//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT64), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AND2_X1   g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(KEYINPUT65), .B1(G567), .B2(new_n454), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n462), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT67), .B1(new_n462), .B2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n479), .A2(KEYINPUT68), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n475), .B1(new_n483), .B2(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g064(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n481), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n463), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n480), .A2(new_n481), .A3(new_n493), .A4(new_n476), .ZN(new_n494));
  INV_X1    g069(.A(G136), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n480), .A2(G2105), .A3(new_n493), .A4(new_n476), .ZN(new_n497));
  OAI221_X1 g072(.A(new_n491), .B1(new_n494), .B2(new_n495), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(G162));
  NAND4_X1  g076(.A1(new_n479), .A2(G126), .A3(G2105), .A4(new_n480), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n481), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT71), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n479), .A2(new_n481), .A3(new_n480), .A4(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n463), .A2(new_n465), .A3(new_n481), .ZN(new_n513));
  INV_X1    g088(.A(G138), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(G164));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(G543), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(G88), .B1(new_n526), .B2(G50), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n526), .A2(G51), .B1(new_n523), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n523), .A2(G89), .A3(new_n524), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g119(.A(KEYINPUT75), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n521), .A2(KEYINPUT5), .A3(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(G543), .B1(new_n521), .B2(KEYINPUT5), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n524), .B(G90), .C1(new_n548), .C2(new_n549), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n524), .A2(G52), .A3(G543), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n554), .A2(KEYINPUT76), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT76), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  AOI22_X1  g134(.A1(new_n525), .A2(G81), .B1(new_n526), .B2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g147(.A1(new_n524), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n573), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n573), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n525), .A2(G91), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n523), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n522), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n577), .B(new_n578), .C1(new_n583), .C2(new_n528), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  NAND2_X1  g161(.A1(new_n525), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n526), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n528), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n523), .A2(new_n524), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n593), .A2(new_n594), .B1(new_n573), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AND2_X1   g173(.A1(new_n523), .A2(G60), .ZN(new_n599));
  AND2_X1   g174(.A1(G72), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n525), .A2(G85), .B1(new_n526), .B2(G47), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n601), .A2(new_n602), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n525), .A2(G92), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n580), .B2(new_n581), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n526), .A2(G54), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n616), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n610), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT81), .B1(new_n624), .B2(G868), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G168), .A2(new_n626), .ZN(new_n627));
  MUX2_X1   g202(.A(new_n625), .B(KEYINPUT81), .S(new_n627), .Z(G297));
  MUX2_X1   g203(.A(new_n625), .B(KEYINPUT81), .S(new_n627), .Z(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n621), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n621), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n481), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n637), .B1(new_n494), .B2(new_n638), .C1(new_n639), .C2(new_n497), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n470), .A2(new_n472), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(KEYINPUT12), .B1(new_n645), .B2(new_n513), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n463), .A2(new_n465), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n647), .A2(new_n648), .A3(new_n481), .A4(new_n644), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT13), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n643), .A2(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n660), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n642), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n689), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n691), .B(new_n694), .C1(new_n686), .C2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT86), .Z(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT85), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n697), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  INV_X1    g284(.A(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT87), .B(G29), .Z(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n481), .A2(G107), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n715), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G119), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n497), .ZN(new_n722));
  INV_X1    g297(.A(G131), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n494), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT89), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n497), .A2(new_n721), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n494), .A2(new_n723), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n720), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n713), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n714), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n711), .B1(new_n712), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n712), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n706), .A2(G22), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G166), .B2(new_n706), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1971), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G1971), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n706), .A2(G6), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n597), .B2(new_n706), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT32), .B(G1981), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n706), .A2(G23), .ZN(new_n743));
  INV_X1    g318(.A(G288), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n706), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT33), .B(G1976), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n737), .A2(new_n738), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT34), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(KEYINPUT34), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n734), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT36), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n706), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n706), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n621), .B2(new_n706), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n706), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n706), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n706), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n706), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(G1966), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n713), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  INV_X1    g347(.A(G140), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n494), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n481), .A2(G116), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n479), .A2(G128), .A3(G2105), .A4(new_n480), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n772), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT91), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n479), .A2(G141), .A3(new_n481), .A4(new_n480), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n479), .A2(G129), .A3(G2105), .A4(new_n480), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT26), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  AOI22_X1  g367(.A1(G105), .A2(new_n473), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT93), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G32), .B(new_n798), .S(G29), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n479), .A2(G139), .A3(new_n481), .A4(new_n480), .ZN(new_n803));
  NAND2_X1  g378(.A1(G115), .A2(G2104), .ZN(new_n804));
  INV_X1    g379(.A(G127), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n466), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G2105), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT25), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n803), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n782), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n782), .B2(G33), .ZN(new_n813));
  INV_X1    g388(.A(G2072), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n566), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G16), .B2(G19), .ZN(new_n818));
  INV_X1    g393(.A(G1341), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G28), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT30), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n821), .B2(KEYINPUT30), .ZN(new_n823));
  OR2_X1    g398(.A1(KEYINPUT31), .A2(G11), .ZN(new_n824));
  NAND2_X1  g399(.A1(KEYINPUT31), .A2(G11), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n819), .A2(new_n818), .B1(new_n813), .B2(new_n814), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n816), .A2(new_n820), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT24), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(G34), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(G34), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n713), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G160), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n782), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G2084), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n641), .B2(new_n713), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n713), .A2(G27), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT96), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G164), .B2(new_n713), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2078), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT97), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n802), .A2(new_n828), .A3(new_n836), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n731), .A2(G35), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G162), .B2(new_n731), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT29), .ZN(new_n845));
  INV_X1    g420(.A(G2090), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n769), .A2(G1966), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT94), .ZN(new_n849));
  AND4_X1   g424(.A1(new_n770), .A2(new_n842), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n752), .A2(new_n763), .A3(new_n850), .ZN(G150));
  INV_X1    g426(.A(G150), .ZN(G311));
  INV_X1    g427(.A(new_n610), .ZN(new_n853));
  INV_X1    g428(.A(new_n620), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT80), .B1(new_n615), .B2(new_n616), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n630), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n525), .A2(G93), .B1(new_n526), .B2(G55), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n528), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n565), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT100), .B(G860), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(new_n516), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n502), .A2(new_n873), .A3(new_n507), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n502), .B2(new_n507), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n781), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n780), .B(new_n872), .C1(new_n874), .C2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n810), .B1(new_n796), .B2(new_n797), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n811), .A2(new_n794), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n479), .A2(G142), .A3(new_n481), .A4(new_n480), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n479), .A2(G130), .A3(G2105), .A4(new_n480), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n888), .A2(new_n481), .A3(G118), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n481), .B2(G118), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n650), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n650), .A2(new_n884), .A3(new_n885), .A4(new_n892), .ZN(new_n896));
  AND4_X1   g471(.A1(new_n725), .A2(new_n729), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n729), .A2(new_n725), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n877), .B(new_n878), .C1(new_n880), .C2(new_n881), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n883), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n833), .B1(new_n499), .B2(new_n500), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n641), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n499), .A2(new_n833), .A3(new_n500), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n883), .A2(new_n900), .ZN(new_n910));
  INV_X1    g485(.A(new_n899), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n883), .A2(new_n899), .A3(new_n900), .A4(KEYINPUT104), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n912), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n907), .A2(new_n908), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT106), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n913), .B(new_n924), .C1(new_n920), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n619), .A2(new_n620), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n624), .B1(new_n929), .B2(new_n853), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n610), .B(G299), .C1(new_n619), .C2(new_n620), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n856), .A2(G299), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n621), .A2(new_n624), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n862), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n632), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n930), .A2(new_n931), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n938), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  NOR2_X1   g517(.A1(G290), .A2(new_n597), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G288), .B1(new_n531), .B2(new_n532), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n531), .A2(new_n532), .A3(G288), .ZN(new_n947));
  AOI21_X1  g522(.A(G305), .B1(new_n605), .B2(new_n606), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n944), .A2(new_n946), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n947), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n951), .A2(new_n945), .B1(new_n943), .B2(new_n948), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n942), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n942), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n861), .A2(new_n626), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n959), .ZN(G331));
  NAND2_X1  g536(.A1(G301), .A2(KEYINPUT108), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n553), .B(new_n963), .C1(new_n556), .C2(new_n557), .ZN(new_n964));
  AND4_X1   g539(.A1(new_n545), .A2(new_n544), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n545), .A2(new_n544), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n937), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(G168), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n544), .A2(new_n962), .A3(new_n545), .A4(new_n964), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n862), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT110), .A3(new_n937), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n969), .A2(new_n940), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n979), .A3(new_n937), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n981), .B2(new_n936), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n953), .B(new_n976), .C1(new_n981), .C2(new_n936), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n979), .B1(new_n974), .B2(new_n937), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT109), .B(new_n862), .C1(new_n971), .C2(new_n972), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n932), .A2(new_n935), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT111), .A3(new_n953), .A4(new_n976), .ZN(new_n991));
  AOI221_X4 g566(.A(G37), .B1(new_n954), .B2(new_n982), .C1(new_n985), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n995));
  AOI21_X1  g570(.A(G37), .B1(new_n985), .B2(new_n991), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n981), .A2(new_n940), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n975), .A2(new_n973), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n936), .B1(new_n998), .B2(new_n969), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n954), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n993), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n994), .B(KEYINPUT44), .C1(new_n995), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n995), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n985), .A2(new_n991), .ZN(new_n1004));
  INV_X1    g579(.A(G37), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n993), .A3(new_n1005), .A4(new_n1000), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n992), .B2(new_n993), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1009));
  OAI22_X1  g584(.A1(new_n1002), .A2(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n876), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G160), .A2(G40), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1996), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT46), .Z(new_n1019));
  XNOR2_X1  g594(.A(new_n780), .B(G2067), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT113), .ZN(new_n1021));
  INV_X1    g596(.A(new_n794), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT123), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT124), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(new_n1024), .A3(KEYINPUT124), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(KEYINPUT47), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n794), .A2(G1996), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1021), .B(new_n1030), .C1(G1996), .C2(new_n798), .ZN(new_n1031));
  INV_X1    g606(.A(new_n712), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n730), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n781), .A2(new_n785), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1017), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n730), .B(new_n1032), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1016), .A2(new_n710), .A3(new_n708), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT125), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT48), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1037), .A2(new_n1016), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1035), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1029), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n597), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n592), .B1(new_n1052), .B2(new_n596), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n596), .A2(new_n1052), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(KEYINPUT116), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1057), .B(new_n1061), .C1(new_n1055), .C2(new_n1058), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1049), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(new_n1065), .A3(new_n1049), .A4(new_n1062), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n744), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1051), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n508), .A2(KEYINPUT101), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n502), .A2(new_n507), .A3(new_n873), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1384), .B1(new_n1073), .B2(new_n872), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1015), .B1(new_n1074), .B2(KEYINPUT45), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1011), .B1(new_n508), .B2(new_n516), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1013), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1971), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1015), .B1(KEYINPUT50), .B2(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n846), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1048), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G303), .A2(G8), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(G166), .B2(new_n1048), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1076), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1015), .B1(new_n1081), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1080), .B1(G2090), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1096), .B2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G286), .A2(new_n1048), .ZN(new_n1099));
  INV_X1    g674(.A(G1966), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1014), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1015), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1013), .B2(new_n1076), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2084), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1082), .A2(new_n1083), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1098), .B(new_n1099), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1091), .B1(new_n1097), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1074), .A2(new_n1102), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(G8), .C1(new_n1068), .C2(G288), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1064), .A2(new_n1066), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1049), .A2(new_n1070), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1117), .B(new_n1099), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT63), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1095), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n846), .A2(new_n1122), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1087), .B(new_n1089), .C1(new_n1123), .C2(new_n1048), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1117), .A2(new_n1124), .A3(new_n1091), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1104), .A2(G168), .A3(new_n1107), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G8), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  AOI21_X1  g704(.A(G168), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1014), .B(new_n1102), .C1(new_n1013), .C2(new_n1076), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1133), .A2(new_n1134), .A3(G2078), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1078), .B2(G2078), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1137));
  INV_X1    g712(.A(G1961), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G171), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1125), .A2(new_n1132), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1129), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1118), .B(new_n1121), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1075), .A2(new_n1077), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1095), .B2(new_n758), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT118), .B(G1956), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(G299), .B(KEYINPUT57), .Z(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1148), .B(new_n1153), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1146), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G1348), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1111), .A2(G2067), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1160), .A2(new_n1161), .A3(KEYINPUT119), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT119), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n856), .B1(new_n1164), .B2(KEYINPUT60), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1166), .B(new_n621), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1165), .A2(new_n1167), .B1(KEYINPUT60), .B2(new_n1164), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT58), .B(G1341), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1078), .A2(G1996), .B1(new_n1047), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n566), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1155), .B1(new_n1164), .B2(new_n856), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1156), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1174), .B2(new_n1156), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1159), .A2(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1134), .A2(G2078), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1075), .A2(new_n1014), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(G301), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1141), .A2(new_n1182), .A3(KEYINPUT122), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1179), .A2(new_n1185), .A3(G301), .A4(new_n1181), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(G171), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1189), .B(KEYINPUT54), .C1(G171), .C2(new_n1140), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1191));
  AND4_X1   g766(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .A4(new_n1125), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1145), .B1(new_n1178), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1037), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G290), .B(new_n710), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1017), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1046), .B1(new_n1193), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g772(.A1(G319), .A2(new_n682), .ZN(new_n1199));
  XNOR2_X1  g773(.A(new_n1199), .B(KEYINPUT126), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n704), .B(new_n1200), .C1(new_n669), .C2(new_n668), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1201), .B1(new_n923), .B2(new_n925), .ZN(new_n1202));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1203));
  INV_X1    g777(.A(new_n1006), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n982), .A2(new_n954), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n993), .B1(new_n996), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g780(.A(new_n1202), .B(new_n1203), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g781(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1203), .B1(new_n1007), .B2(new_n1202), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n1208), .A2(new_n1209), .ZN(G308));
  OAI21_X1  g784(.A(new_n1202), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1211), .A2(KEYINPUT127), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(new_n1207), .ZN(G225));
endmodule


