//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT64), .A2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT64), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR3_X1   g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G143), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n193), .A2(new_n194), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n202), .A2(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT3), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT3), .A2(G107), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(G104), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT82), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT82), .A2(G104), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G101), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n213), .B2(new_n219), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n219), .A3(new_n223), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT4), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n210), .B(new_n222), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT10), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(G128), .B1(new_n204), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n196), .B2(new_n201), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT64), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT64), .A2(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(G143), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n200), .A3(new_n199), .A4(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n223), .B1(G104), .B2(G107), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n228), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT64), .B(G146), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n204), .B1(new_n246), .B2(new_n195), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n237), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT10), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n227), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n252), .A2(G134), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(G134), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n251), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n254), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n256), .B2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n251), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n250), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n255), .A2(new_n251), .A3(new_n260), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n227), .A2(new_n243), .A3(new_n270), .A4(new_n249), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT81), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n244), .A2(new_n248), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n242), .B1(new_n237), .B2(new_n231), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n267), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n270), .B2(KEYINPUT83), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n242), .B(new_n237), .C1(new_n247), .C2(new_n245), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n242), .B2(new_n238), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n284), .B1(new_n288), .B2(new_n267), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n271), .B(new_n277), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n279), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n192), .B1(new_n291), .B2(new_n190), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n268), .A2(new_n271), .A3(new_n277), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n285), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n267), .A3(new_n284), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n227), .A2(new_n243), .A3(new_n249), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n270), .ZN(new_n297));
  OAI211_X1 g111(.A(G469), .B(new_n293), .C1(new_n297), .C2(new_n277), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n189), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(KEYINPUT70), .A2(G237), .ZN(new_n300));
  NOR2_X1   g114(.A1(KEYINPUT70), .A2(G237), .ZN(new_n301));
  OAI211_X1 g115(.A(G214), .B(new_n273), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n195), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT70), .B(G237), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n304), .A2(G143), .A3(G214), .A4(new_n273), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT18), .A2(G131), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n198), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n317), .A2(new_n246), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT76), .B1(new_n206), .B2(new_n310), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT89), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n309), .A2(new_n321), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT70), .A2(G237), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT70), .A2(G237), .ZN(new_n332));
  AOI21_X1  g146(.A(G953), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(G143), .B1(new_n333), .B2(G214), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n302), .A2(new_n195), .ZN(new_n335));
  OAI21_X1  g149(.A(G131), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n303), .A2(new_n305), .A3(new_n251), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n306), .A2(KEYINPUT17), .A3(G131), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n317), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n198), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n310), .B2(KEYINPUT16), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n341), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n198), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT90), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n339), .A2(new_n340), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n327), .A2(new_n330), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n330), .B1(new_n327), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n191), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G475), .ZN(new_n357));
  NOR2_X1   g171(.A1(G475), .A2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n317), .B(KEYINPUT19), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n246), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n346), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n336), .A2(new_n338), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n318), .B1(new_n317), .B2(new_n246), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n206), .A2(new_n310), .A3(KEYINPUT76), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n311), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n325), .B1(new_n369), .B2(new_n309), .ZN(new_n370));
  INV_X1    g184(.A(new_n326), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n330), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n353), .B(new_n330), .C1(new_n370), .C2(new_n371), .ZN(new_n375));
  AOI211_X1 g189(.A(KEYINPUT20), .B(new_n359), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n324), .A2(new_n326), .B1(new_n363), .B2(new_n362), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n375), .B1(new_n330), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n379), .B2(new_n358), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n357), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT73), .B(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(new_n187), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n235), .B2(G143), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n195), .A2(KEYINPUT91), .A3(G128), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n235), .A2(G143), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT92), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT92), .B1(new_n387), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n256), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(KEYINPUT13), .A3(new_n386), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G134), .ZN(new_n397));
  XNOR2_X1  g211(.A(G116), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(G107), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n396), .B2(G134), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n392), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G116), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n216), .B1(new_n408), .B2(KEYINPUT14), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n398), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n388), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(G134), .A3(new_n389), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n392), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n383), .B1(new_n406), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n383), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n419), .B(new_n416), .C1(new_n403), .C2(new_n405), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n191), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n392), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT93), .B1(new_n404), .B2(new_n392), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n419), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n406), .A2(new_n417), .A3(new_n383), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n423), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n381), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n299), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  INV_X1    g253(.A(G116), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(KEYINPUT2), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n438), .A2(new_n443), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n244), .A2(new_n436), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n242), .B2(KEYINPUT86), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT8), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G119), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G116), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n444), .B(new_n446), .C1(new_n441), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n447), .A2(new_n437), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(new_n222), .C1(new_n226), .C2(new_n224), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n442), .A2(new_n455), .A3(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(G116), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(G119), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(G113), .B(new_n461), .C1(new_n464), .C2(new_n442), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n225), .A2(new_n465), .A3(new_n458), .A4(new_n241), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT84), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n448), .A2(new_n468), .A3(new_n225), .A4(new_n241), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n460), .A2(new_n467), .A3(new_n452), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n234), .A2(new_n200), .A3(new_n199), .A4(new_n203), .ZN(new_n471));
  INV_X1    g285(.A(new_n209), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n247), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n273), .A2(G224), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT7), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n315), .B(new_n237), .C1(new_n245), .C2(new_n247), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n454), .B(new_n470), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT87), .B1(new_n480), .B2(new_n191), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(KEYINPUT87), .A3(new_n191), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n485));
  INV_X1    g299(.A(new_n452), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n470), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n485), .B(new_n486), .C1(KEYINPUT85), .C2(new_n488), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n474), .A2(new_n477), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n273), .A2(G224), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n484), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n481), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n483), .B(KEYINPUT88), .Z(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(G234), .A2(G237), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(G952), .A3(new_n273), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(G902), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT21), .B(G898), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G214), .B1(G237), .B2(G902), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n501), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n435), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G472), .A2(G902), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n254), .B2(new_n257), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n266), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n248), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n207), .A2(new_n209), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n471), .B(new_n518), .C1(new_n269), .C2(new_n261), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT68), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT68), .B1(new_n457), .B2(new_n458), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT69), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n517), .A2(new_n519), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n519), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n459), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT28), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n267), .A2(new_n210), .B1(new_n516), .B2(new_n248), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT28), .B1(new_n531), .B2(new_n522), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n333), .A2(G210), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT27), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n514), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n532), .B1(new_n529), .B2(KEYINPUT28), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n541), .A2(KEYINPUT71), .A3(new_n538), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n544));
  OR2_X1    g358(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n517), .A2(new_n519), .A3(new_n545), .A4(new_n544), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n459), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n524), .A2(new_n526), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n551), .A3(new_n538), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT31), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n527), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n554), .A2(new_n547), .B1(new_n457), .B2(new_n458), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n550), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n538), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT32), .B(new_n513), .C1(new_n543), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n539), .B1(new_n541), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n524), .B(new_n526), .C1(new_n531), .C2(new_n522), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n532), .B1(new_n563), .B2(KEYINPUT28), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n555), .A2(new_n550), .A3(new_n538), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n566), .B2(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  INV_X1    g383(.A(new_n513), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n553), .A2(new_n558), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n534), .A2(new_n514), .A3(new_n539), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT71), .B1(new_n541), .B2(new_n538), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n570), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n576));
  OAI211_X1 g390(.A(new_n560), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n382), .B1(G234), .B2(new_n191), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n455), .B2(G128), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n455), .B2(G128), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n235), .A2(G119), .ZN(new_n584));
  NOR2_X1   g398(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n581), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G110), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT24), .B(G110), .Z(new_n588));
  XNOR2_X1  g402(.A(G119), .B(G128), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n587), .B(new_n590), .C1(new_n346), .C2(new_n348), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT22), .B(G137), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT75), .B(G110), .Z(new_n595));
  OAI22_X1  g409(.A1(new_n586), .A2(new_n595), .B1(new_n589), .B2(new_n588), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n366), .A2(new_n367), .ZN(new_n597));
  AND4_X1   g411(.A1(KEYINPUT77), .A2(new_n596), .A3(new_n597), .A4(new_n351), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n366), .A2(new_n367), .B1(new_n347), .B2(G146), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT77), .B1(new_n599), .B2(new_n596), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n591), .B(new_n594), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n587), .A2(new_n590), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n351), .B2(new_n350), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(new_n597), .A3(new_n351), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(KEYINPUT77), .A3(new_n596), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n594), .B(KEYINPUT78), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n601), .B(new_n191), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT25), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n579), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT25), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n578), .A2(G902), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n601), .B(new_n617), .C1(new_n608), .C2(new_n609), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n577), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(KEYINPUT80), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT80), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n577), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n512), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  OAI21_X1  g439(.A(new_n191), .B1(new_n543), .B2(new_n559), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n575), .B1(new_n626), .B2(G472), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n627), .A2(new_n619), .A3(new_n299), .ZN(new_n628));
  INV_X1    g442(.A(new_n510), .ZN(new_n629));
  INV_X1    g443(.A(new_n483), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n497), .B2(new_n481), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n631), .B2(new_n496), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n509), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n422), .A2(new_n191), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n430), .B2(new_n422), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT33), .B1(new_n418), .B2(new_n420), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n428), .A2(new_n429), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(G478), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n381), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n628), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AOI22_X1  g459(.A1(new_n424), .A2(new_n432), .B1(G475), .B2(new_n356), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n379), .A2(new_n358), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n379), .A2(new_n377), .A3(new_n358), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(KEYINPUT94), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT94), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n380), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n646), .A2(new_n650), .A3(new_n509), .A4(new_n652), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n632), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n628), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  AND2_X1   g474(.A1(new_n501), .A2(new_n510), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT36), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n609), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n608), .B(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n614), .A2(new_n615), .B1(new_n664), .B2(new_n617), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n665), .A2(new_n381), .A3(new_n433), .A4(new_n508), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n627), .A2(new_n661), .A3(new_n299), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NAND2_X1  g483(.A1(new_n664), .A2(new_n617), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n616), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n271), .A2(new_n277), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n295), .B2(new_n294), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n277), .B1(new_n268), .B2(new_n271), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n190), .B(new_n191), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n192), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n298), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n188), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n503), .B(KEYINPUT96), .Z(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(G900), .B2(new_n505), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n646), .A2(new_n650), .A3(new_n652), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n631), .A2(new_n496), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n510), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n577), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XNOR2_X1  g500(.A(new_n680), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n299), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT40), .Z(new_n689));
  INV_X1    g503(.A(KEYINPUT98), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n575), .A2(new_n576), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n556), .A2(new_n539), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n191), .B1(new_n563), .B2(new_n538), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n692), .A2(KEYINPUT97), .A3(new_n560), .A4(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n560), .B(new_n695), .C1(new_n575), .C2(new_n576), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT97), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n689), .A2(new_n690), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n501), .B(KEYINPUT38), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n381), .A2(new_n433), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n510), .A2(new_n702), .A3(new_n665), .A4(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n691), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NAND4_X1  g520(.A1(new_n381), .A2(new_n639), .A3(new_n635), .A4(new_n680), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n678), .A2(new_n707), .A3(new_n683), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n577), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT99), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n577), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NOR2_X1   g528(.A1(new_n291), .A2(new_n190), .ZN(new_n715));
  INV_X1    g529(.A(new_n675), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n189), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n577), .A2(new_n619), .A3(new_n642), .A4(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n718), .B(new_n720), .ZN(G15));
  NAND3_X1  g535(.A1(new_n577), .A2(new_n619), .A3(new_n717), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n656), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n440), .ZN(G18));
  NOR2_X1   g538(.A1(new_n715), .A2(new_n716), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n188), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n683), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n577), .A2(new_n666), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NOR2_X1   g543(.A1(new_n564), .A2(new_n538), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n513), .B1(new_n559), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n571), .B2(new_n574), .ZN(new_n732));
  INV_X1    g546(.A(G472), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n619), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n717), .A2(new_n703), .A3(new_n509), .A4(new_n632), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT101), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT101), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  OAI211_X1 g554(.A(new_n671), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n707), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n727), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  AOI22_X1  g559(.A1(new_n575), .A2(KEYINPUT32), .B1(G472), .B2(new_n568), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n575), .B2(KEYINPUT32), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n513), .B1(new_n543), .B2(new_n559), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT32), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n298), .A2(KEYINPUT102), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n271), .B1(new_n286), .B2(new_n289), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n278), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n756), .A3(G469), .A4(new_n293), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n753), .A2(new_n675), .A3(new_n757), .A4(new_n676), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n189), .B1(new_n758), .B2(KEYINPUT103), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n510), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n292), .A2(new_n762), .A3(new_n757), .A4(new_n753), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n707), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n752), .A2(new_n764), .A3(new_n619), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n764), .A2(new_n577), .A3(new_n619), .A4(new_n743), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n761), .A2(new_n766), .A3(new_n763), .A4(new_n759), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(KEYINPUT106), .A3(new_n619), .A4(new_n752), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  XNOR2_X1  g590(.A(new_n681), .B(KEYINPUT107), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n764), .A3(new_n577), .A4(new_n619), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  AND2_X1   g593(.A1(new_n755), .A2(new_n293), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n780), .B2(KEYINPUT45), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n784), .B2(new_n676), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n716), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n676), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n189), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(new_n687), .A3(new_n761), .ZN(new_n789));
  INV_X1    g603(.A(new_n640), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n790), .A2(KEYINPUT43), .A3(new_n381), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT43), .B1(new_n790), .B2(new_n381), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n671), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n793), .A2(new_n794), .A3(new_n627), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n793), .B2(new_n627), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n789), .A2(new_n795), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT109), .B(G137), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G39));
  NAND2_X1  g616(.A1(new_n786), .A2(new_n787), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n188), .ZN(new_n804));
  AND2_X1   g618(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n788), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n577), .A2(new_n619), .A3(new_n707), .A4(new_n760), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  XOR2_X1   g627(.A(new_n725), .B(KEYINPUT49), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n619), .A2(new_n510), .A3(new_n188), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n381), .A3(new_n790), .ZN(new_n816));
  OR4_X1    g630(.A1(new_n700), .A2(new_n702), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n577), .A2(new_n708), .A3(new_n711), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n711), .B1(new_n577), .B2(new_n708), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n685), .B(new_n744), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n680), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n671), .A2(KEYINPUT112), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n665), .B2(new_n680), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n703), .A2(new_n632), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n829), .A3(new_n763), .A4(new_n759), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n696), .B2(new_n699), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n819), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n830), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n700), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n744), .A2(new_n685), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n713), .A4(KEYINPUT52), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT101), .ZN(new_n838));
  INV_X1    g652(.A(new_n734), .ZN(new_n839));
  INV_X1    g653(.A(new_n735), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n841), .A2(new_n736), .B1(new_n722), .B2(new_n656), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n424), .A2(new_n432), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(new_n381), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n511), .B1(new_n844), .B2(new_n641), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n627), .A3(new_n619), .A4(new_n299), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n718), .A2(new_n846), .A3(new_n667), .A4(new_n728), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n764), .A2(new_n742), .A3(new_n743), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n823), .B1(new_n356), .B2(G475), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n843), .A2(new_n650), .A3(new_n652), .A4(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n678), .A2(new_n851), .A3(new_n760), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(new_n577), .A3(KEYINPUT111), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT111), .B1(new_n852), .B2(new_n577), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n778), .B(new_n849), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n848), .A2(new_n856), .A3(new_n775), .A4(new_n624), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n818), .B1(new_n837), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n832), .A2(new_n836), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n667), .A2(new_n718), .A3(new_n846), .A4(new_n728), .ZN(new_n861));
  INV_X1    g675(.A(new_n723), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n624), .A2(new_n861), .A3(new_n862), .A4(new_n739), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n855), .B1(new_n864), .B2(new_n774), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n863), .A3(KEYINPUT53), .A4(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n858), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n859), .B1(new_n858), .B2(new_n866), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n856), .A2(new_n775), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n861), .A2(new_n624), .A3(new_n862), .A4(new_n739), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n873), .B2(new_n860), .ZN(new_n874));
  AND4_X1   g688(.A1(KEYINPUT53), .A2(new_n860), .A3(new_n863), .A4(new_n865), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n858), .A2(new_n859), .A3(new_n866), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT113), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n679), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n791), .A2(new_n880), .A3(new_n792), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n734), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n715), .A2(new_n716), .A3(new_n188), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n761), .B(new_n882), .C1(new_n810), .C2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n702), .A2(new_n510), .A3(new_n726), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT50), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(KEYINPUT50), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n726), .A2(new_n760), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n887), .A2(new_n888), .B1(new_n742), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n619), .A3(new_n504), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n700), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n640), .A2(new_n381), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n884), .A2(new_n892), .A3(KEYINPUT51), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n752), .A2(new_n619), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT115), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT115), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT48), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n273), .A2(G952), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n700), .A2(new_n641), .A3(new_n893), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n907), .B(new_n908), .C1(new_n727), .C2(new_n882), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n897), .A2(new_n904), .A3(new_n906), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n804), .A2(new_n805), .ZN(new_n913));
  INV_X1    g727(.A(new_n809), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n883), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n882), .A2(new_n761), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n896), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n892), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n911), .B(new_n912), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT114), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n910), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n879), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n817), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n273), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n191), .B1(new_n858), .B2(new_n866), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n490), .A2(new_n491), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n494), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n928), .A2(new_n936), .A3(new_n499), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n928), .B2(new_n499), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(new_n192), .B(KEYINPUT57), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n876), .B2(new_n877), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n858), .A2(new_n859), .A3(new_n866), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n945), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n673), .A2(new_n674), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n928), .A2(new_n783), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n926), .B1(new_n953), .B2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n374), .A3(new_n375), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .A4(new_n379), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n927), .A3(new_n958), .ZN(G60));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n636), .A2(new_n638), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n634), .B(KEYINPUT59), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT119), .B1(new_n867), .B2(new_n868), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n948), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n926), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n946), .B2(new_n949), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n927), .ZN(new_n970));
  INV_X1    g784(.A(new_n963), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n870), .B2(new_n878), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n962), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(new_n858), .A2(new_n866), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT122), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n975), .A2(new_n981), .A3(new_n664), .A4(new_n977), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n980), .A2(new_n927), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n975), .A2(new_n664), .A3(new_n977), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT122), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n986), .ZN(new_n991));
  INV_X1    g805(.A(new_n988), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n990), .B(new_n991), .C1(new_n983), .C2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n989), .A2(new_n993), .ZN(G66));
  INV_X1    g808(.A(new_n507), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n273), .B1(new_n995), .B2(G224), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n872), .B2(new_n273), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n930), .B1(G898), .B2(new_n273), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(G69));
  NOR2_X1   g813(.A1(new_n546), .A2(new_n548), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT124), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(new_n360), .Z(new_n1002));
  OAI211_X1 g816(.A(G900), .B(G953), .C1(new_n1002), .C2(G227), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G227), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n844), .A2(new_n641), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT125), .Z(new_n1006));
  NOR2_X1   g820(.A1(new_n688), .A2(new_n760), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1006), .B(new_n1007), .C1(new_n621), .C2(new_n623), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n800), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  INV_X1    g824(.A(new_n822), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n705), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT62), .Z(new_n1013));
  NAND3_X1  g827(.A1(new_n1010), .A2(new_n812), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1002), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n788), .A2(new_n687), .A3(new_n898), .A4(new_n829), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n812), .A2(new_n778), .A3(new_n1017), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n775), .A2(new_n1018), .A3(new_n800), .A4(new_n1011), .ZN(new_n1019));
  AOI21_X1  g833(.A(G953), .B1(new_n1019), .B2(new_n1002), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1004), .B1(new_n1016), .B2(new_n1020), .ZN(G72));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n566), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1010), .A2(new_n693), .A3(new_n812), .A4(new_n1013), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n872), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n693), .A2(new_n566), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AOI211_X1 g842(.A(new_n1025), .B(new_n1028), .C1(new_n858), .C2(new_n866), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1027), .B(KEYINPUT127), .Z(new_n1030));
  AND2_X1   g844(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NOR4_X1   g845(.A1(new_n1024), .A2(new_n926), .A3(new_n1029), .A4(new_n1031), .ZN(G57));
endmodule


