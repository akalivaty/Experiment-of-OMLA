//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT83), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(KEYINPUT22), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  AND2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT24), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n218), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n218), .A2(new_n224), .A3(new_n229), .A4(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n221), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT65), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n236), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT64), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n226), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G183gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n255), .A3(new_n226), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(KEYINPUT28), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n245), .B(new_n228), .C1(new_n252), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n234), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n215), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(KEYINPUT72), .B(new_n261), .C1(new_n234), .C2(new_n259), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n226), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n256), .A2(new_n257), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n245), .A4(new_n228), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n234), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n216), .B1(new_n267), .B2(new_n268), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n270), .B1(new_n273), .B2(new_n245), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n261), .B(KEYINPUT71), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n214), .B1(new_n265), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n272), .B2(new_n274), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n273), .A2(new_n245), .B1(new_n232), .B2(new_n233), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n261), .B1(new_n281), .B2(KEYINPUT29), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n282), .A3(new_n214), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT37), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n207), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n214), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n281), .B2(new_n261), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n260), .A2(new_n215), .A3(new_n262), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n234), .A3(new_n271), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n276), .B1(new_n291), .B2(new_n266), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n286), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n293), .A2(KEYINPUT83), .A3(KEYINPUT37), .A4(new_n283), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT38), .B1(new_n285), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n214), .C1(new_n289), .C2(new_n292), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n286), .B1(new_n265), .B2(new_n278), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n282), .A3(new_n286), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT73), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT37), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n301), .A2(KEYINPUT84), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT84), .B1(new_n301), .B2(new_n302), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n206), .B(new_n295), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT0), .ZN(new_n308));
  XNOR2_X1  g107(.A(G57gat), .B(G85gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT67), .B(G113gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n315), .B(new_n323), .C1(new_n324), .C2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n328));
  OAI21_X1  g127(.A(G162gat), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n330));
  OR2_X1    g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G155gat), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336));
  AND4_X1   g135(.A1(new_n331), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n338), .A3(new_n336), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n335), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n330), .A2(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n326), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(G155gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n338), .B1(new_n345), .B2(G162gat), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n342), .B(new_n344), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n312), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n348), .A4(new_n326), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n351), .B2(new_n326), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n323), .A2(new_n315), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n361));
  OAI21_X1  g160(.A(G120gat), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n359), .A2(new_n362), .B1(new_n316), .B2(new_n321), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n341), .A3(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n350), .B2(new_n353), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n355), .A4(new_n356), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n356), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n351), .B(new_n326), .ZN(new_n374));
  INV_X1    g173(.A(new_n356), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n355), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n306), .B(new_n311), .C1(new_n372), .C2(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n368), .A2(new_n371), .B1(new_n373), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT82), .B1(new_n379), .B2(new_n310), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT6), .B1(new_n379), .B2(new_n310), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n379), .A2(new_n310), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT6), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n301), .A2(new_n385), .A3(new_n205), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n301), .B2(new_n205), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n305), .A2(new_n382), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT38), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n301), .A2(new_n302), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n301), .A2(KEYINPUT84), .A3(new_n302), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n205), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n301), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT37), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n342), .B1(new_n214), .B2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n351), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n214), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n403), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n407), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n406), .B1(KEYINPUT80), .B2(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n206), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n301), .A2(KEYINPUT30), .A3(new_n205), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n388), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n363), .B1(KEYINPUT3), .B2(new_n351), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT77), .B1(new_n424), .B2(new_n348), .ZN(new_n425));
  INV_X1    g224(.A(new_n353), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n366), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT81), .B1(new_n427), .B2(new_n375), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n369), .A2(new_n429), .A3(new_n356), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(KEYINPUT81), .A3(new_n375), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n369), .B2(new_n356), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n374), .A2(new_n375), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT39), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n310), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n431), .A2(new_n435), .A3(KEYINPUT40), .A4(new_n310), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n380), .A4(new_n378), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n417), .B1(new_n422), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n202), .B1(new_n399), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n305), .A2(new_n388), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n382), .A2(new_n384), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n206), .B(new_n397), .C1(new_n303), .C2(new_n304), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT38), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n413), .A2(new_n416), .ZN(new_n448));
  INV_X1    g247(.A(new_n440), .ZN(new_n449));
  INV_X1    g248(.A(new_n420), .ZN(new_n450));
  INV_X1    g249(.A(new_n387), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n301), .A2(new_n385), .A3(new_n205), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n421), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n448), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n455), .A3(KEYINPUT85), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n457));
  INV_X1    g256(.A(new_n381), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n384), .B1(new_n458), .B2(new_n383), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n459), .A3(new_n460), .A4(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n448), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n290), .A2(new_n363), .A3(new_n234), .A4(new_n271), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n291), .A2(new_n326), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n271), .A2(new_n234), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n363), .A4(new_n290), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n471), .A3(new_n465), .ZN(new_n473));
  INV_X1    g272(.A(new_n468), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT34), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT33), .B1(new_n473), .B2(new_n474), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI211_X1 g284(.A(new_n477), .B(new_n485), .C1(new_n473), .C2(new_n474), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n476), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n473), .A2(new_n474), .ZN(new_n488));
  INV_X1    g287(.A(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT32), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n475), .A3(new_n472), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT69), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n476), .A2(new_n486), .ZN(new_n494));
  INV_X1    g293(.A(new_n478), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(new_n482), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT69), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n487), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n498), .A2(new_n490), .B1(new_n475), .B2(new_n472), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n492), .B1(new_n483), .B2(new_n491), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n494), .A2(KEYINPUT69), .A3(new_n498), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT70), .B1(new_n507), .B2(KEYINPUT36), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n498), .B2(new_n494), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT36), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n442), .A2(new_n456), .A3(new_n462), .A4(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n500), .A2(new_n454), .A3(new_n448), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n417), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n461), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(new_n334), .ZN(new_n521));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  INV_X1    g324(.A(G64gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G57gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(G57gat), .ZN(new_n528));
  INV_X1    g327(.A(G57gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT93), .A3(G64gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G71gat), .B(G78gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(KEYINPUT95), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n536), .B1(KEYINPUT9), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT96), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n554));
  OR3_X1    g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G127gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n559));
  AND2_X1   g358(.A1(KEYINPUT90), .A2(G1gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(KEYINPUT90), .A2(G1gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT16), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT91), .ZN(new_n563));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G1gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n565), .A2(G8gat), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(G8gat), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n319), .A3(new_n556), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n558), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n558), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n524), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n573), .A3(new_n523), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT87), .B(G29gat), .Z(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(KEYINPUT88), .A3(G36gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT87), .B(G29gat), .ZN(new_n583));
  INV_X1    g382(.A(G36gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(G29gat), .A2(G36gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT14), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n590));
  INV_X1    g389(.A(G43gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n592));
  XOR2_X1   g391(.A(G43gat), .B(G50gat), .Z(new_n593));
  OAI211_X1 g392(.A(new_n590), .B(new_n592), .C1(new_n593), .C2(KEYINPUT89), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n596), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT8), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n602), .B(new_n604), .C1(G85gat), .C2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n600), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(new_n599), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT92), .B1(new_n610), .B2(KEYINPUT17), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n598), .C2(new_n599), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(new_n607), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n609), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n625), .A2(KEYINPUT98), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n609), .B(new_n620), .C1(new_n615), .C2(new_n618), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(KEYINPUT98), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT99), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n622), .A2(new_n626), .A3(new_n627), .A4(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n607), .B1(new_n549), .B2(new_n551), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n548), .A2(new_n607), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n552), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT100), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(KEYINPUT101), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n645), .B(new_n651), .C1(KEYINPUT101), .C2(new_n650), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n579), .A2(new_n635), .A3(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n570), .B(new_n616), .C1(new_n611), .C2(new_n614), .ZN(new_n658));
  NAND2_X1  g457(.A1(G229gat), .A2(G233gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n600), .A2(new_n568), .A3(new_n569), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n658), .A2(KEYINPUT18), .A3(new_n659), .A4(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n570), .A2(new_n610), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n660), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n659), .B(KEYINPUT13), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G169gat), .B(G197gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT12), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n663), .A2(new_n664), .A3(new_n668), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n661), .A2(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n678), .B2(new_n664), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n657), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n519), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n459), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n566), .ZN(G1324gat));
  INV_X1    g483(.A(G8gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n682), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n454), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n682), .A2(new_n422), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n689), .ZN(G1325gat));
  AOI21_X1  g490(.A(G15gat), .B1(new_n686), .B2(new_n507), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT102), .ZN(new_n693));
  INV_X1    g492(.A(new_n511), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n686), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n417), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n519), .A2(new_n634), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n635), .B1(new_n512), .B2(new_n518), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n579), .A2(new_n680), .A3(new_n655), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n580), .B1(new_n708), .B2(new_n459), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n704), .A2(new_n707), .ZN(new_n710));
  INV_X1    g509(.A(new_n459), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n583), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1328gat));
  OAI21_X1  g513(.A(G36gat), .B1(new_n708), .B2(new_n422), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n584), .A3(new_n454), .ZN(new_n716));
  AND2_X1   g515(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n715), .B(new_n719), .C1(new_n717), .C2(new_n716), .ZN(G1329gat));
  NAND2_X1  g519(.A1(new_n694), .A2(G43gat), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n710), .A2(new_n507), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n708), .A2(new_n721), .B1(G43gat), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n708), .B2(new_n417), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n417), .A2(G50gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  AOI21_X1  g532(.A(new_n634), .B1(new_n578), .B2(new_n576), .ZN(new_n734));
  AND4_X1   g533(.A1(new_n519), .A2(new_n680), .A3(new_n734), .A4(new_n655), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n711), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n454), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT49), .B(G64gat), .Z(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n735), .A2(new_n694), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n500), .A2(G71gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(G71gat), .B1(new_n735), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n735), .A2(new_n448), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT106), .B(G78gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  INV_X1    g547(.A(G85gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n711), .A2(new_n749), .A3(new_n655), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n519), .A2(KEYINPUT107), .A3(new_n634), .ZN(new_n752));
  INV_X1    g551(.A(new_n680), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n579), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n759));
  INV_X1    g558(.A(new_n754), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n704), .B2(KEYINPUT107), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n751), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n761), .A3(KEYINPUT51), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n750), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n760), .A2(new_n656), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n706), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n749), .B1(new_n769), .B2(new_n711), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT109), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n750), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n765), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT108), .B1(new_n764), .B2(new_n765), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n706), .A2(new_n768), .ZN(new_n777));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777), .B2(new_n459), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n771), .A2(new_n779), .ZN(G1336gat));
  NOR2_X1   g579(.A1(new_n422), .A2(G92gat), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n655), .B(new_n781), .C1(new_n758), .C2(new_n762), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n703), .A2(new_n454), .A3(new_n705), .A4(new_n768), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g585(.A1(new_n500), .A2(G99gat), .A3(new_n656), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n773), .B2(new_n774), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n777), .B2(new_n511), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NOR2_X1   g589(.A1(new_n417), .A2(G106gat), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n655), .B(new_n791), .C1(new_n758), .C2(new_n762), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n703), .A2(new_n448), .A3(new_n705), .A4(new_n768), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g595(.A1(new_n657), .A2(new_n753), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n639), .A2(new_n643), .A3(new_n640), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n645), .A2(new_n799), .A3(KEYINPUT54), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n648), .B1(new_n653), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(new_n652), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n666), .A2(new_n667), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n673), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n676), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n800), .A2(new_n802), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n634), .A2(new_n804), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n655), .A2(new_n676), .A3(new_n807), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n677), .B2(new_n679), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n803), .A2(new_n652), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n635), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n798), .B1(new_n817), .B2(new_n579), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n711), .ZN(new_n819));
  INV_X1    g618(.A(new_n516), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n422), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n324), .A3(new_n753), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n513), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n680), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n314), .A3(new_n655), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n824), .B2(new_n656), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT110), .ZN(G1341gat));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n319), .A3(new_n579), .ZN(new_n831));
  INV_X1    g630(.A(new_n579), .ZN(new_n832));
  OAI21_X1  g631(.A(G127gat), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1342gat));
  NOR2_X1   g633(.A1(new_n635), .A2(new_n454), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n821), .A2(new_n317), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT56), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n513), .A3(new_n634), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n836), .A2(KEYINPUT56), .B1(new_n840), .B2(G134gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1343gat));
  INV_X1    g641(.A(G141gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n511), .A2(new_n711), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n454), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n800), .B2(new_n802), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n663), .A2(new_n664), .A3(new_n668), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n674), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n676), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n850), .A2(new_n804), .B1(new_n655), .B2(new_n808), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n634), .B1(new_n851), .B2(KEYINPUT113), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n816), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n812), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n798), .B1(new_n855), .B2(new_n579), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .A3(new_n448), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n818), .A2(new_n448), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n846), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n843), .B1(new_n861), .B2(new_n753), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n844), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n680), .A2(G141gat), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n863), .A2(new_n422), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT58), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n863), .B(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n422), .A3(new_n864), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n866), .B1(new_n871), .B2(new_n862), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n656), .A2(G148gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n422), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  INV_X1    g674(.A(new_n859), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n816), .A2(new_n635), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n804), .A2(new_n808), .A3(new_n634), .A4(new_n811), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n579), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n448), .B(new_n876), .C1(new_n879), .C2(new_n797), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n818), .A2(new_n882), .A3(new_n448), .A4(new_n876), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n657), .B2(new_n753), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n734), .A2(KEYINPUT116), .A3(new_n680), .A4(new_n656), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n855), .B2(new_n579), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n448), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n655), .B(new_n845), .C1(new_n884), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n875), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n875), .A2(G148gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n861), .B2(new_n655), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n874), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n874), .B(new_n897), .C1(new_n892), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1345gat));
  NOR2_X1   g698(.A1(new_n832), .A2(new_n345), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n868), .A2(new_n422), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n861), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n345), .B1(new_n902), .B2(new_n832), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1346gat));
  NAND3_X1  g703(.A1(new_n868), .A2(new_n332), .A3(new_n835), .ZN(new_n905));
  OAI21_X1  g704(.A(G162gat), .B1(new_n902), .B2(new_n635), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  NAND3_X1  g706(.A1(new_n507), .A2(new_n454), .A3(new_n459), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT120), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n448), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n818), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n220), .A3(new_n680), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n818), .A2(new_n459), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n516), .A2(new_n422), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT118), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n753), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n918), .B2(new_n220), .ZN(G1348gat));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n221), .A3(new_n655), .ZN(new_n920));
  OAI21_X1  g719(.A(G176gat), .B1(new_n911), .B2(new_n656), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n579), .A2(new_n251), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n818), .A2(new_n459), .A3(new_n915), .A4(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n911), .B2(new_n832), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n818), .A2(KEYINPUT122), .A3(new_n579), .A4(new_n910), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(G183gat), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n923), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n923), .A3(new_n930), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n932), .A2(new_n933), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(new_n933), .ZN(new_n935));
  NAND2_X1  g734(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(new_n931), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n934), .A2(new_n937), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n226), .A3(new_n634), .ZN(new_n939));
  OAI21_X1  g738(.A(G190gat), .B1(new_n911), .B2(new_n635), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1351gat));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n511), .A2(new_n448), .A3(new_n454), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n818), .B(new_n459), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n753), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n884), .A2(new_n890), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n511), .A2(new_n459), .A3(new_n454), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT127), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n753), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n949), .B1(new_n947), .B2(new_n954), .ZN(G1352gat));
  NAND3_X1  g754(.A1(new_n950), .A2(new_n655), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n946), .A2(new_n958), .A3(new_n655), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n209), .A3(new_n579), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n950), .A2(new_n579), .A3(new_n952), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NAND3_X1  g766(.A1(new_n946), .A2(new_n210), .A3(new_n634), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n634), .A3(new_n952), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(new_n210), .ZN(G1355gat));
endmodule


