//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(KEYINPUT85), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(new_n208), .B2(new_n209), .ZN(new_n216));
  AOI211_X1 g015(.A(KEYINPUT86), .B(new_n206), .C1(new_n212), .C2(new_n213), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n204), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n210), .B(KEYINPUT88), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n204), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(KEYINPUT15), .B2(new_n203), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n219), .A2(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(KEYINPUT89), .A3(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n225), .A2(new_n226), .ZN(new_n232));
  NAND2_X1  g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT7), .ZN(new_n234));
  INV_X1    g033(.A(G99gat), .ZN(new_n235));
  INV_X1    g034(.A(G106gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT8), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT95), .B(G92gat), .Z(new_n238));
  OAI211_X1 g037(.A(new_n234), .B(new_n237), .C1(G85gat), .C2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G99gat), .B(G106gat), .Z(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  NOR2_X1   g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT41), .ZN(new_n245));
  INV_X1    g044(.A(new_n225), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n239), .B(new_n240), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G190gat), .B(G218gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT96), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n244), .A2(KEYINPUT41), .ZN(new_n253));
  XNOR2_X1  g052(.A(G134gat), .B(G162gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT97), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n251), .ZN(new_n258));
  INV_X1    g057(.A(new_n243), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n248), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n255), .A2(KEYINPUT97), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G71gat), .A2(G78gat), .ZN(new_n267));
  OR2_X1    g066(.A1(G71gat), .A2(G78gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT9), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271));
  INV_X1    g070(.A(G64gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(G57gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(G57gat), .B2(new_n272), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(G57gat), .B2(new_n272), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n267), .B(new_n268), .C1(new_n277), .C2(new_n269), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT93), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G127gat), .ZN(new_n285));
  XOR2_X1   g084(.A(G183gat), .B(G211gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT16), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G1gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(G1gat), .B2(new_n288), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(G8gat), .Z(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n280), .B2(new_n281), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT94), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n294), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n287), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT93), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n279), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n247), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n241), .A2(new_n279), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT10), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT10), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n280), .A2(new_n247), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G230gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n307), .A2(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G176gat), .B(G204gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT100), .ZN(new_n317));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n314), .A3(new_n321), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n323), .A2(KEYINPUT101), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT101), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n266), .A2(new_n302), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G197gat), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT11), .B(G169gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  NOR2_X1   g133(.A1(new_n246), .A2(new_n292), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n292), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT91), .B1(new_n225), .B2(new_n337), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n225), .A2(KEYINPUT91), .A3(new_n337), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT90), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT13), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n232), .A2(new_n337), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n342), .B(new_n335), .C1(new_n231), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n346), .B2(KEYINPUT18), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n231), .A2(new_n345), .ZN(new_n348));
  INV_X1    g147(.A(new_n342), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n349), .A4(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n334), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n336), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT18), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n334), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n350), .A4(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n329), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n361));
  OR2_X1    g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT27), .B(G183gat), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT28), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G183gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT27), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G183gat), .ZN(new_n379));
  AND4_X1   g178(.A1(KEYINPUT28), .A2(new_n377), .A3(new_n379), .A4(new_n374), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n372), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT69), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n385), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n381), .A2(new_n391), .A3(KEYINPUT70), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n379), .A3(new_n374), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT28), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n373), .A2(KEYINPUT28), .A3(new_n374), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n396), .A2(new_n397), .B1(G183gat), .B2(G190gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n385), .A2(new_n387), .A3(new_n390), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G169gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT65), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT65), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G169gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT23), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT66), .B(G176gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT67), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT68), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n388), .B2(KEYINPUT23), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(KEYINPUT68), .C1(G169gat), .C2(G176gat), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n410), .A2(new_n412), .B1(G169gat), .B2(G176gat), .ZN(new_n413));
  AND2_X1   g212(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT65), .B(G169gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT67), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(KEYINPUT23), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n372), .ZN(new_n421));
  NAND3_X1  g220(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n408), .A2(new_n413), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n412), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n427), .A2(new_n423), .A3(new_n383), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n388), .B2(KEYINPUT23), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n401), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(KEYINPUT29), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n424), .A2(new_n425), .B1(new_n428), .B2(new_n430), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n381), .A2(new_n391), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n371), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT70), .B1(new_n381), .B2(new_n391), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n398), .A2(new_n393), .A3(new_n399), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n443), .B2(new_n436), .ZN(new_n444));
  INV_X1    g243(.A(new_n437), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n432), .A2(new_n445), .A3(new_n433), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n371), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND4_X1  g249(.A1(new_n440), .A2(new_n447), .A3(KEYINPUT30), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  INV_X1    g251(.A(new_n447), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n439), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n447), .A3(new_n450), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G141gat), .B(G148gat), .Z(new_n461));
  INV_X1    g260(.A(KEYINPUT2), .ZN(new_n462));
  INV_X1    g261(.A(G162gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G155gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n296), .A2(G162gat), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n461), .A2(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G120gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G113gat), .ZN(new_n469));
  INV_X1    g268(.A(G113gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G120gat), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT1), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(G127gat), .A2(G134gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(G127gat), .A2(G134gat), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT1), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n476), .A2(KEYINPUT71), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n473), .A2(new_n474), .B1(KEYINPUT71), .B2(new_n476), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n469), .A2(new_n471), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT1), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(G148gat), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G141gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(G148gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(KEYINPUT75), .A2(G162gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT2), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n491), .A2(new_n464), .A3(new_n465), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n489), .A2(KEYINPUT76), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT76), .B1(new_n489), .B2(new_n492), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n467), .B(new_n482), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n498));
  AND2_X1   g297(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n487), .B1(new_n501), .B2(G148gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n491), .A2(new_n464), .A3(new_n465), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT76), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n466), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n507));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n497), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT77), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n482), .B1(new_n506), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n467), .B1(new_n493), .B2(new_n494), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n509), .A2(new_n516), .A3(KEYINPUT80), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n507), .A3(new_n508), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n508), .ZN(new_n527));
  INV_X1    g326(.A(new_n495), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n505), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n482), .B1(new_n529), .B2(new_n467), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT79), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT79), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(new_n527), .C1(new_n528), .C2(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n516), .A3(KEYINPUT78), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n526), .A2(new_n535), .A3(KEYINPUT5), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT0), .ZN(new_n539));
  XNOR2_X1  g338(.A(G57gat), .B(G85gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n522), .B2(new_n537), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n537), .ZN(new_n547));
  INV_X1    g346(.A(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT6), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n460), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(G50gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n370), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n506), .B1(new_n556), .B2(new_n511), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n506), .A2(new_n511), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n370), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n554), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n557), .A2(new_n559), .A3(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(G228gat), .A2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G22gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n561), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n561), .B2(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G227gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(new_n311), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n482), .B1(new_n443), .B2(new_n436), .ZN(new_n573));
  INV_X1    g372(.A(new_n482), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n432), .A2(new_n574), .A3(new_n441), .A4(new_n442), .ZN(new_n575));
  AOI211_X1 g374(.A(KEYINPUT34), .B(new_n572), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n572), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n401), .B2(new_n432), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n443), .A2(new_n436), .A3(new_n482), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT34), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n575), .A3(new_n572), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585));
  XOR2_X1   g384(.A(G15gat), .B(G43gat), .Z(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G99gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n584), .B(KEYINPUT32), .C1(new_n585), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(KEYINPUT32), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n585), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n580), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n583), .A2(new_n590), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(new_n576), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT34), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n570), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n551), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n547), .A2(new_n548), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n543), .A3(new_n542), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n549), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n609));
  AND4_X1   g408(.A1(new_n570), .A2(new_n595), .A3(new_n602), .A4(new_n609), .ZN(new_n610));
  AND4_X1   g409(.A1(KEYINPUT84), .A2(new_n608), .A3(new_n460), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n459), .B1(new_n607), .B2(new_n549), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT84), .B1(new_n612), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n605), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n570), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n545), .B1(new_n458), .B2(new_n455), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n497), .A2(new_n507), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n508), .B1(new_n617), .B2(new_n516), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n514), .A2(new_n574), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n508), .A3(new_n495), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT39), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT82), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT82), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n625), .A3(KEYINPUT39), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n620), .B(new_n541), .C1(new_n627), .C2(new_n618), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT40), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n615), .B1(new_n616), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT37), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n454), .B1(new_n632), .B2(new_n450), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n443), .A2(new_n436), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n432), .A2(new_n445), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n634), .A2(new_n433), .B1(new_n635), .B2(new_n435), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n447), .B1(new_n636), .B2(new_n371), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT37), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n631), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n452), .B1(new_n637), .B2(KEYINPUT37), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n444), .A2(new_n370), .A3(new_n446), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n641), .B(KEYINPUT37), .C1(new_n636), .C2(new_n370), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n456), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n607), .A3(new_n549), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n595), .A2(new_n602), .A3(KEYINPUT36), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648));
  INV_X1    g447(.A(new_n595), .ZN(new_n649));
  INV_X1    g448(.A(new_n602), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n630), .A2(new_n646), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n551), .A2(new_n615), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n614), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n360), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n608), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n459), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(G8gat), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n662), .A2(new_n661), .A3(new_n665), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  NOR2_X1   g468(.A1(new_n649), .A2(new_n650), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n657), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n647), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT103), .Z(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n657), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n656), .A2(new_n570), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  AOI21_X1  g478(.A(new_n266), .B1(new_n614), .B2(new_n654), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n359), .A2(new_n302), .A3(new_n327), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n208), .A3(new_n658), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n263), .A2(new_n265), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n551), .A2(new_n688), .A3(new_n615), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n612), .B2(new_n570), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n652), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n614), .B2(new_n691), .ZN(new_n692));
  OAI22_X1  g491(.A1(KEYINPUT105), .A2(new_n692), .B1(new_n680), .B2(new_n686), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(KEYINPUT105), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n681), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT106), .B(new_n681), .C1(new_n693), .C2(new_n694), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n700), .A3(new_n608), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n685), .B1(new_n701), .B2(new_n208), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n682), .A2(G36gat), .A3(new_n460), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n698), .A2(new_n700), .A3(new_n460), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n209), .ZN(G1329gat));
  OAI21_X1  g505(.A(G43gat), .B1(new_n695), .B2(new_n672), .ZN(new_n707));
  INV_X1    g506(.A(new_n670), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n682), .A2(G43gat), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n673), .A3(new_n699), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n695), .B2(new_n570), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n682), .A2(G50gat), .A3(new_n570), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n615), .A3(new_n699), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(G50gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g521(.A1(new_n359), .A2(new_n266), .A3(new_n302), .A4(new_n327), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n614), .B2(new_n691), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n658), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g525(.A(new_n460), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT107), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n670), .B(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(G71gat), .B1(new_n724), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n673), .A2(G71gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n724), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n724), .A2(new_n615), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g539(.A1(new_n693), .A2(new_n694), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n358), .A2(new_n302), .A3(new_n328), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743), .B2(new_n608), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n614), .A2(new_n691), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n266), .A2(new_n358), .A3(new_n302), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n745), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n608), .A2(G85gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n327), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n755), .ZN(G1336gat));
  OAI211_X1 g555(.A(new_n459), .B(new_n742), .C1(new_n693), .C2(new_n694), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n238), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n460), .A2(G92gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n752), .A2(new_n327), .A3(new_n753), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n327), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n764), .A3(new_n750), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n745), .B(new_n746), .C1(KEYINPUT111), .C2(KEYINPUT51), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n769), .B2(KEYINPUT52), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n757), .B2(new_n238), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n759), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n762), .B1(new_n770), .B2(new_n773), .ZN(G1337gat));
  NOR3_X1   g573(.A1(new_n743), .A2(new_n235), .A3(new_n672), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n752), .A2(new_n670), .A3(new_n327), .A4(new_n753), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n235), .B2(new_n776), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n741), .A2(new_n615), .A3(new_n742), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G106gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n328), .A2(G106gat), .A3(new_n570), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n752), .A2(new_n753), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n766), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n778), .A2(G106gat), .B1(new_n784), .B2(new_n781), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n780), .B2(new_n785), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n305), .A2(new_n306), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n309), .B1(new_n787), .B2(new_n308), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n313), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n321), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n313), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(KEYINPUT54), .A3(new_n312), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n324), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n352), .B2(new_n357), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n349), .B1(new_n348), .B2(new_n336), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n340), .A2(new_n343), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n333), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n357), .A2(new_n327), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n266), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n257), .A2(new_n264), .A3(new_n260), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n264), .B1(new_n257), .B2(new_n260), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n801), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n811), .A2(new_n357), .A3(new_n812), .A4(new_n805), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n302), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n329), .A2(new_n358), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n658), .A2(new_n460), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n604), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n358), .A2(new_n470), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n820), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n359), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n822), .A2(new_n823), .B1(new_n826), .B2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n824), .B2(new_n328), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n327), .A2(new_n468), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n822), .B2(new_n830), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832));
  INV_X1    g631(.A(new_n302), .ZN(new_n833));
  OR4_X1    g632(.A1(KEYINPUT116), .A2(new_n824), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n821), .A2(new_n302), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n835), .B2(new_n832), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n832), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(G1342gat));
  NAND3_X1  g637(.A1(new_n818), .A2(new_n811), .A3(new_n820), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n839), .A2(G134gat), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g639(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n839), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT117), .B1(new_n839), .B2(G134gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n839), .A2(G134gat), .ZN(new_n845));
  OAI221_X1 g644(.A(new_n842), .B1(new_n843), .B2(new_n844), .C1(new_n845), .C2(new_n841), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n819), .A2(new_n673), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n615), .B(new_n847), .C1(new_n814), .C2(new_n816), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n358), .A2(new_n486), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT119), .Z(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n795), .A2(new_n797), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n352), .B2(new_n357), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n266), .B1(new_n854), .B2(new_n807), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n813), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n816), .B1(new_n856), .B2(new_n833), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n857), .B2(new_n570), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n615), .C1(new_n814), .C2(new_n816), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n858), .A2(new_n358), .A3(new_n860), .A4(new_n847), .ZN(new_n861));
  INV_X1    g660(.A(new_n501), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n851), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n864), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n851), .B(new_n866), .C1(new_n861), .C2(new_n862), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  OR3_X1    g667(.A1(new_n848), .A2(G148gat), .A3(new_n328), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n615), .B1(new_n814), .B2(new_n816), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n358), .A2(new_n852), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n811), .B1(new_n872), .B2(new_n806), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n357), .A2(new_n805), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n266), .A2(new_n801), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n833), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n817), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n570), .A2(KEYINPUT57), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n871), .A2(KEYINPUT57), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n327), .A3(new_n847), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n870), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n870), .A2(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n858), .A2(new_n860), .A3(new_n847), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n327), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n869), .B1(new_n881), .B2(new_n885), .ZN(G1345gat));
  OAI21_X1  g685(.A(G155gat), .B1(new_n883), .B2(new_n833), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n302), .A2(new_n296), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n848), .B2(new_n888), .ZN(G1346gat));
  XNOR2_X1  g688(.A(KEYINPUT75), .B(G162gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n883), .B2(new_n266), .ZN(new_n891));
  OR4_X1    g690(.A1(new_n673), .A2(new_n266), .A3(new_n819), .A4(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n871), .B2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n658), .A2(new_n460), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n733), .A2(new_n570), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n818), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n359), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n604), .A2(new_n460), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n608), .B(new_n898), .C1(new_n814), .C2(new_n816), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n417), .A3(new_n358), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT121), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n896), .A2(new_n416), .A3(new_n328), .ZN(new_n904));
  AOI21_X1  g703(.A(G176gat), .B1(new_n900), .B2(new_n327), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1349gat));
  NAND2_X1  g705(.A1(new_n302), .A2(new_n373), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n900), .A2(KEYINPUT122), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n899), .B2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G183gat), .B1(new_n896), .B2(new_n833), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n374), .A3(new_n811), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n811), .B(new_n895), .C1(new_n814), .C2(new_n816), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G190gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT123), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(G190gat), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n922), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n919), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  AOI21_X1  g727(.A(new_n658), .B1(new_n815), .B2(new_n817), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n673), .A2(new_n460), .A3(new_n570), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n931), .A2(G197gat), .A3(new_n359), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n877), .A2(new_n878), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n894), .A2(new_n672), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT124), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n937), .B2(new_n359), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n359), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n328), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n931), .A2(KEYINPUT62), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n937), .B2(new_n328), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT62), .B1(new_n931), .B2(new_n943), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1353gat));
  NOR2_X1   g746(.A1(new_n935), .A2(new_n833), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n879), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(KEYINPUT126), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT63), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n949), .B(new_n952), .C1(KEYINPUT126), .C2(new_n951), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n929), .A2(new_n950), .A3(new_n302), .A4(new_n930), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1354gat));
  NOR2_X1   g757(.A1(new_n931), .A2(new_n266), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n811), .A2(G218gat), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n959), .A2(G218gat), .B1(new_n937), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(G1355gat));
endmodule


