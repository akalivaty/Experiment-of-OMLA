

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n537), .A2(G2104), .ZN(n889) );
  NOR2_X1 U556 ( .A1(n593), .A2(n552), .ZN(n797) );
  BUF_X1 U557 ( .A(n723), .Z(n724) );
  AND2_X2 U558 ( .A1(n535), .A2(G2105), .ZN(n885) );
  XNOR2_X1 U559 ( .A(n620), .B(KEYINPUT28), .ZN(n650) );
  XNOR2_X1 U560 ( .A(n539), .B(n538), .ZN(n541) );
  AND2_X1 U561 ( .A1(n625), .A2(G1996), .ZN(n624) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT99), .ZN(n667) );
  NAND2_X1 U563 ( .A1(n665), .A2(n664), .ZN(n688) );
  NAND2_X1 U564 ( .A1(n659), .A2(n658), .ZN(n660) );
  AND2_X1 U565 ( .A1(n702), .A2(n701), .ZN(n703) );
  INV_X1 U566 ( .A(G2105), .ZN(n537) );
  AND2_X1 U567 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X2 U568 ( .A1(n721), .A2(n616), .ZN(n625) );
  AND2_X1 U569 ( .A1(n763), .A2(n753), .ZN(n523) );
  AND2_X1 U570 ( .A1(n719), .A2(n526), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT66), .B(n536), .Z(n525) );
  OR2_X1 U572 ( .A1(n701), .A2(n718), .ZN(n526) );
  XNOR2_X1 U573 ( .A(KEYINPUT14), .B(n626), .ZN(n527) );
  AND2_X1 U574 ( .A1(n802), .A2(G43), .ZN(n528) );
  AND2_X1 U575 ( .A1(G137), .A2(n723), .ZN(n529) );
  XOR2_X1 U576 ( .A(KEYINPUT31), .B(n672), .Z(n530) );
  XOR2_X1 U577 ( .A(n668), .B(n667), .Z(n531) );
  INV_X1 U578 ( .A(n950), .ZN(n633) );
  AND2_X1 U579 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U580 ( .A1(n636), .A2(n635), .ZN(n637) );
  INV_X1 U581 ( .A(KEYINPUT98), .ZN(n654) );
  XNOR2_X1 U582 ( .A(n660), .B(KEYINPUT29), .ZN(n665) );
  INV_X1 U583 ( .A(n625), .ZN(n681) );
  XNOR2_X1 U584 ( .A(n700), .B(KEYINPUT101), .ZN(n702) );
  NAND2_X1 U585 ( .A1(n681), .A2(G8), .ZN(n680) );
  NAND2_X1 U586 ( .A1(n885), .A2(G125), .ZN(n536) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n538) );
  INV_X1 U588 ( .A(KEYINPUT68), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n532), .B(KEYINPUT17), .ZN(n533) );
  NAND2_X1 U590 ( .A1(G160), .A2(G40), .ZN(n721) );
  XNOR2_X1 U591 ( .A(n534), .B(n533), .ZN(n723) );
  INV_X1 U592 ( .A(G2104), .ZN(n535) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n553), .Z(n805) );
  NOR2_X1 U594 ( .A1(G651), .A2(n593), .ZN(n802) );
  NOR2_X1 U595 ( .A1(n631), .A2(n528), .ZN(n632) );
  NAND2_X1 U596 ( .A1(n548), .A2(n547), .ZN(G160) );
  NAND2_X1 U597 ( .A1(n527), .A2(n632), .ZN(n950) );
  NOR2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n529), .A2(n525), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G101), .A2(n889), .ZN(n539) );
  AND2_X1 U601 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U602 ( .A1(G113), .A2(n886), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n546) );
  INV_X1 U604 ( .A(n546), .ZN(n545) );
  INV_X1 U605 ( .A(KEYINPUT65), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n546), .A2(KEYINPUT65), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT0), .B(G543), .Z(n593) );
  INV_X1 U609 ( .A(G651), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G78), .A2(n797), .ZN(n550) );
  NOR2_X1 U611 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U612 ( .A1(G91), .A2(n798), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U614 ( .A(KEYINPUT71), .B(n551), .ZN(n557) );
  NOR2_X1 U615 ( .A1(G543), .A2(n552), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G65), .A2(n805), .ZN(n555) );
  NAND2_X1 U617 ( .A1(G53), .A2(n802), .ZN(n554) );
  AND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U620 ( .A1(G126), .A2(n885), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G114), .A2(n886), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G138), .A2(n723), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n889), .A2(G102), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U626 ( .A(KEYINPUT93), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n564) );
  NOR2_X1 U628 ( .A1(n565), .A2(n564), .ZN(G164) );
  NAND2_X1 U629 ( .A1(G64), .A2(n805), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G52), .A2(n802), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G77), .A2(n797), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G90), .A2(n798), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(n571), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(G171) );
  NAND2_X1 U638 ( .A1(G63), .A2(n805), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G51), .A2(n802), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT6), .B(n576), .ZN(n584) );
  NAND2_X1 U642 ( .A1(G89), .A2(n798), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G76), .A2(n797), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT5), .B(n582), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT7), .B(n585), .Z(G168) );
  NAND2_X1 U651 ( .A1(G75), .A2(n797), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G88), .A2(n798), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G62), .A2(n805), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G50), .A2(n802), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(G166) );
  INV_X1 U658 ( .A(G166), .ZN(G303) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(n592) );
  XNOR2_X1 U660 ( .A(KEYINPUT76), .B(n592), .ZN(G286) );
  NAND2_X1 U661 ( .A1(n593), .A2(G87), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G49), .A2(n802), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G74), .A2(G651), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U665 ( .A1(n805), .A2(n596), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U667 ( .A(KEYINPUT83), .B(n599), .Z(G288) );
  NAND2_X1 U668 ( .A1(G61), .A2(n805), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G86), .A2(n798), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U671 ( .A(KEYINPUT84), .B(n602), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n797), .A2(G73), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT2), .B(n603), .Z(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n802), .A2(G48), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(G305) );
  NAND2_X1 U677 ( .A1(G60), .A2(n805), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G47), .A2(n802), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G72), .A2(n797), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT69), .B(n610), .ZN(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n798), .A2(G85), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(G290) );
  INV_X1 U685 ( .A(G299), .ZN(n937) );
  NOR2_X1 U686 ( .A1(G164), .A2(G1384), .ZN(n722) );
  INV_X1 U687 ( .A(n722), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n625), .A2(G2072), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT27), .ZN(n619) );
  INV_X1 U690 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U691 ( .A1(n969), .A2(n625), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n937), .A2(n621), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n937), .A2(n621), .ZN(n622) );
  OR2_X1 U695 ( .A1(n650), .A2(n622), .ZN(n659) );
  INV_X1 U696 ( .A(KEYINPUT26), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n636) );
  NAND2_X1 U698 ( .A1(n681), .A2(G1341), .ZN(n634) );
  NAND2_X1 U699 ( .A1(G56), .A2(n805), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n798), .A2(G81), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G68), .A2(n797), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U704 ( .A(KEYINPUT13), .B(n630), .Z(n631) );
  XNOR2_X1 U705 ( .A(n637), .B(KEYINPUT64), .ZN(n653) );
  NAND2_X1 U706 ( .A1(G66), .A2(n805), .ZN(n639) );
  NAND2_X1 U707 ( .A1(G92), .A2(n798), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U709 ( .A1(G79), .A2(n797), .ZN(n641) );
  NAND2_X1 U710 ( .A1(G54), .A2(n802), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(n949) );
  NAND2_X1 U715 ( .A1(n653), .A2(n949), .ZN(n649) );
  NOR2_X1 U716 ( .A1(n625), .A2(G1348), .ZN(n647) );
  NOR2_X1 U717 ( .A1(G2067), .A2(n681), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n652) );
  INV_X1 U720 ( .A(n650), .ZN(n651) );
  AND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n653), .A2(n949), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n625), .A2(G1961), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n661), .B(KEYINPUT97), .ZN(n663) );
  XNOR2_X1 U727 ( .A(G2078), .B(KEYINPUT25), .ZN(n987) );
  NAND2_X1 U728 ( .A1(n625), .A2(n987), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U730 ( .A1(n669), .A2(G171), .ZN(n664) );
  NOR2_X1 U731 ( .A1(G1966), .A2(n680), .ZN(n675) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n681), .ZN(n677) );
  NOR2_X1 U733 ( .A1(n675), .A2(n677), .ZN(n666) );
  NAND2_X1 U734 ( .A1(G8), .A2(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(G168), .A2(n531), .ZN(n671) );
  NOR2_X1 U736 ( .A1(G171), .A2(n669), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n688), .A2(n530), .ZN(n674) );
  INV_X1 U739 ( .A(KEYINPUT100), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n679) );
  NAND2_X1 U742 ( .A1(G8), .A2(n677), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n696) );
  INV_X1 U744 ( .A(G8), .ZN(n686) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n680), .ZN(n683) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n681), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n684), .A2(G303), .ZN(n685) );
  OR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n689) );
  AND2_X1 U750 ( .A1(n530), .A2(n689), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n693) );
  INV_X1 U752 ( .A(n689), .ZN(n691) );
  AND2_X1 U753 ( .A1(G286), .A2(G8), .ZN(n690) );
  OR2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n694), .B(KEYINPUT32), .ZN(n695) );
  NAND2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n715) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n942) );
  NOR2_X1 U759 ( .A1(G1971), .A2(G303), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n942), .A2(n697), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n715), .A2(n698), .ZN(n699) );
  NAND2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NAND2_X1 U763 ( .A1(n699), .A2(n943), .ZN(n700) );
  INV_X1 U764 ( .A(n680), .ZN(n701) );
  NOR2_X1 U765 ( .A1(KEYINPUT33), .A2(n703), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n704), .B(KEYINPUT102), .ZN(n705) );
  XNOR2_X1 U767 ( .A(G1981), .B(G305), .ZN(n935) );
  NOR2_X1 U768 ( .A1(n705), .A2(n935), .ZN(n709) );
  NAND2_X1 U769 ( .A1(n942), .A2(KEYINPUT33), .ZN(n706) );
  XNOR2_X1 U770 ( .A(KEYINPUT103), .B(n706), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n707), .A2(n701), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n720) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT24), .ZN(n711) );
  NAND2_X1 U775 ( .A1(n711), .A2(n701), .ZN(n719) );
  NOR2_X1 U776 ( .A1(G2090), .A2(G303), .ZN(n712) );
  XNOR2_X1 U777 ( .A(KEYINPUT104), .B(n712), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n713), .A2(G8), .ZN(n714) );
  XOR2_X1 U779 ( .A(KEYINPUT105), .B(n714), .Z(n716) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U781 ( .A(KEYINPUT106), .B(n717), .Z(n718) );
  NAND2_X1 U782 ( .A1(n720), .A2(n524), .ZN(n754) );
  NOR2_X1 U783 ( .A1(n722), .A2(n721), .ZN(n766) );
  NAND2_X1 U784 ( .A1(n889), .A2(G104), .ZN(n726) );
  NAND2_X1 U785 ( .A1(G140), .A2(n724), .ZN(n725) );
  NAND2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n727), .ZN(n732) );
  NAND2_X1 U788 ( .A1(G128), .A2(n885), .ZN(n729) );
  NAND2_X1 U789 ( .A1(G116), .A2(n886), .ZN(n728) );
  NAND2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U791 ( .A(KEYINPUT35), .B(n730), .Z(n731) );
  NOR2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U793 ( .A(KEYINPUT36), .B(n733), .ZN(n909) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(G2067), .ZN(n755) );
  NOR2_X1 U795 ( .A1(n909), .A2(n755), .ZN(n1010) );
  NAND2_X1 U796 ( .A1(n766), .A2(n1010), .ZN(n763) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(KEYINPUT95), .Z(n735) );
  NAND2_X1 U798 ( .A1(G105), .A2(n889), .ZN(n734) );
  XNOR2_X1 U799 ( .A(n735), .B(n734), .ZN(n742) );
  NAND2_X1 U800 ( .A1(n885), .A2(G129), .ZN(n737) );
  NAND2_X1 U801 ( .A1(G141), .A2(n724), .ZN(n736) );
  NAND2_X1 U802 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U803 ( .A1(n886), .A2(G117), .ZN(n738) );
  XOR2_X1 U804 ( .A(KEYINPUT94), .B(n738), .Z(n739) );
  NOR2_X1 U805 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U806 ( .A1(n742), .A2(n741), .ZN(n900) );
  NAND2_X1 U807 ( .A1(G1996), .A2(n900), .ZN(n743) );
  XOR2_X1 U808 ( .A(KEYINPUT96), .B(n743), .Z(n751) );
  NAND2_X1 U809 ( .A1(n889), .A2(G95), .ZN(n745) );
  NAND2_X1 U810 ( .A1(G131), .A2(n724), .ZN(n744) );
  NAND2_X1 U811 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U812 ( .A1(G119), .A2(n885), .ZN(n747) );
  NAND2_X1 U813 ( .A1(G107), .A2(n886), .ZN(n746) );
  NAND2_X1 U814 ( .A1(n747), .A2(n746), .ZN(n748) );
  OR2_X1 U815 ( .A1(n749), .A2(n748), .ZN(n904) );
  AND2_X1 U816 ( .A1(n904), .A2(G1991), .ZN(n750) );
  NOR2_X1 U817 ( .A1(n751), .A2(n750), .ZN(n758) );
  XOR2_X1 U818 ( .A(G1986), .B(G290), .Z(n953) );
  NAND2_X1 U819 ( .A1(n758), .A2(n953), .ZN(n752) );
  NAND2_X1 U820 ( .A1(n752), .A2(n766), .ZN(n753) );
  NAND2_X1 U821 ( .A1(n754), .A2(n523), .ZN(n769) );
  NAND2_X1 U822 ( .A1(n909), .A2(n755), .ZN(n1009) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n900), .ZN(n756) );
  XOR2_X1 U824 ( .A(KEYINPUT107), .B(n756), .Z(n1025) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n904), .ZN(n1013) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n757) );
  NOR2_X1 U827 ( .A1(n1013), .A2(n757), .ZN(n759) );
  INV_X1 U828 ( .A(n758), .ZN(n1017) );
  NOR2_X1 U829 ( .A1(n759), .A2(n1017), .ZN(n760) );
  NOR2_X1 U830 ( .A1(n1025), .A2(n760), .ZN(n761) );
  XNOR2_X1 U831 ( .A(KEYINPUT39), .B(n761), .ZN(n762) );
  XNOR2_X1 U832 ( .A(n762), .B(KEYINPUT108), .ZN(n764) );
  NAND2_X1 U833 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U834 ( .A1(n1009), .A2(n765), .ZN(n767) );
  NAND2_X1 U835 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U836 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U837 ( .A(n770), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U841 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U842 ( .A(G223), .ZN(n843) );
  NAND2_X1 U843 ( .A1(n843), .A2(G567), .ZN(n772) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n778) );
  OR2_X1 U846 ( .A1(n950), .A2(n778), .ZN(G153) );
  INV_X1 U847 ( .A(G171), .ZN(G301) );
  NAND2_X1 U848 ( .A1(G301), .A2(G868), .ZN(n773) );
  XNOR2_X1 U849 ( .A(n773), .B(KEYINPUT72), .ZN(n775) );
  OR2_X1 U850 ( .A1(G868), .A2(n949), .ZN(n774) );
  NAND2_X1 U851 ( .A1(n775), .A2(n774), .ZN(G284) );
  NAND2_X1 U852 ( .A1(G868), .A2(G286), .ZN(n777) );
  INV_X1 U853 ( .A(G868), .ZN(n821) );
  NAND2_X1 U854 ( .A1(G299), .A2(n821), .ZN(n776) );
  NAND2_X1 U855 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n778), .A2(G559), .ZN(n779) );
  NAND2_X1 U857 ( .A1(n779), .A2(n949), .ZN(n780) );
  XNOR2_X1 U858 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U859 ( .A1(G868), .A2(n950), .ZN(n781) );
  XOR2_X1 U860 ( .A(KEYINPUT77), .B(n781), .Z(n784) );
  NAND2_X1 U861 ( .A1(G868), .A2(n949), .ZN(n782) );
  NOR2_X1 U862 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U863 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U864 ( .A(KEYINPUT78), .B(n785), .ZN(G282) );
  XOR2_X1 U865 ( .A(G2100), .B(KEYINPUT80), .Z(n795) );
  NAND2_X1 U866 ( .A1(G99), .A2(n889), .ZN(n787) );
  NAND2_X1 U867 ( .A1(G111), .A2(n886), .ZN(n786) );
  NAND2_X1 U868 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U869 ( .A1(n885), .A2(G123), .ZN(n788) );
  XOR2_X1 U870 ( .A(KEYINPUT18), .B(n788), .Z(n789) );
  NOR2_X1 U871 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U872 ( .A1(G135), .A2(n724), .ZN(n791) );
  NAND2_X1 U873 ( .A1(n792), .A2(n791), .ZN(n1014) );
  XNOR2_X1 U874 ( .A(KEYINPUT79), .B(n1014), .ZN(n793) );
  XNOR2_X1 U875 ( .A(n793), .B(G2096), .ZN(n794) );
  NAND2_X1 U876 ( .A1(n795), .A2(n794), .ZN(G156) );
  NAND2_X1 U877 ( .A1(n949), .A2(G559), .ZN(n819) );
  XNOR2_X1 U878 ( .A(n950), .B(n819), .ZN(n796) );
  NOR2_X1 U879 ( .A1(n796), .A2(G860), .ZN(n809) );
  NAND2_X1 U880 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U881 ( .A1(G93), .A2(n798), .ZN(n799) );
  NAND2_X1 U882 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U883 ( .A(n801), .B(KEYINPUT81), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G55), .A2(n802), .ZN(n803) );
  NAND2_X1 U885 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U886 ( .A1(n805), .A2(G67), .ZN(n806) );
  XOR2_X1 U887 ( .A(KEYINPUT82), .B(n806), .Z(n807) );
  OR2_X1 U888 ( .A1(n808), .A2(n807), .ZN(n822) );
  XOR2_X1 U889 ( .A(n809), .B(n822), .Z(G145) );
  XOR2_X1 U890 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n811) );
  XNOR2_X1 U891 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n810) );
  XNOR2_X1 U892 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U893 ( .A(G166), .B(n812), .ZN(n814) );
  XNOR2_X1 U894 ( .A(n950), .B(n937), .ZN(n813) );
  XNOR2_X1 U895 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U896 ( .A(n822), .B(n815), .ZN(n816) );
  XNOR2_X1 U897 ( .A(G305), .B(n816), .ZN(n817) );
  XNOR2_X1 U898 ( .A(n817), .B(G290), .ZN(n818) );
  XNOR2_X1 U899 ( .A(n818), .B(G288), .ZN(n912) );
  XNOR2_X1 U900 ( .A(n912), .B(n819), .ZN(n820) );
  NOR2_X1 U901 ( .A1(n821), .A2(n820), .ZN(n824) );
  NOR2_X1 U902 ( .A1(G868), .A2(n822), .ZN(n823) );
  NOR2_X1 U903 ( .A1(n824), .A2(n823), .ZN(G295) );
  XNOR2_X1 U904 ( .A(KEYINPUT20), .B(KEYINPUT89), .ZN(n827) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n825) );
  XNOR2_X1 U906 ( .A(n825), .B(KEYINPUT88), .ZN(n826) );
  XNOR2_X1 U907 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n828), .ZN(n829) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U910 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U912 ( .A1(G132), .A2(G82), .ZN(n831) );
  XNOR2_X1 U913 ( .A(n831), .B(KEYINPUT22), .ZN(n832) );
  XNOR2_X1 U914 ( .A(n832), .B(KEYINPUT90), .ZN(n833) );
  NOR2_X1 U915 ( .A1(G218), .A2(n833), .ZN(n834) );
  NAND2_X1 U916 ( .A1(G96), .A2(n834), .ZN(n849) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n849), .ZN(n835) );
  XNOR2_X1 U918 ( .A(KEYINPUT91), .B(n835), .ZN(n840) );
  NAND2_X1 U919 ( .A1(G69), .A2(G120), .ZN(n836) );
  NOR2_X1 U920 ( .A1(G237), .A2(n836), .ZN(n837) );
  NAND2_X1 U921 ( .A1(G108), .A2(n837), .ZN(n848) );
  NAND2_X1 U922 ( .A1(G567), .A2(n848), .ZN(n838) );
  XOR2_X1 U923 ( .A(KEYINPUT92), .B(n838), .Z(n839) );
  NOR2_X1 U924 ( .A1(n840), .A2(n839), .ZN(G319) );
  INV_X1 U925 ( .A(G319), .ZN(n842) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U927 ( .A1(n842), .A2(n841), .ZN(n847) );
  NAND2_X1 U928 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U931 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n845) );
  XOR2_X1 U933 ( .A(KEYINPUT111), .B(n845), .Z(n846) );
  NAND2_X1 U934 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U936 ( .A(G132), .ZN(G219) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G82), .ZN(G220) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2678), .B(KEYINPUT42), .Z(n851) );
  XNOR2_X1 U943 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U944 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U945 ( .A(KEYINPUT112), .B(G2090), .Z(n853) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U948 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U949 ( .A(G2100), .B(G2096), .ZN(n856) );
  XNOR2_X1 U950 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U951 ( .A(G2084), .B(G2078), .Z(n858) );
  XNOR2_X1 U952 ( .A(n859), .B(n858), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1976), .B(G1981), .Z(n861) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1956), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U956 ( .A(n862), .B(G2474), .Z(n864) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U959 ( .A(KEYINPUT41), .B(G1971), .Z(n866) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1961), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U962 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G124), .A2(n885), .ZN(n869) );
  XNOR2_X1 U964 ( .A(n869), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G100), .A2(n889), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n870), .B(KEYINPUT114), .ZN(n871) );
  NAND2_X1 U967 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U968 ( .A1(n886), .A2(G112), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G136), .A2(n724), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U971 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U972 ( .A1(n889), .A2(G103), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G139), .A2(n724), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U975 ( .A1(n885), .A2(G127), .ZN(n879) );
  XOR2_X1 U976 ( .A(KEYINPUT115), .B(n879), .Z(n881) );
  NAND2_X1 U977 ( .A1(n886), .A2(G115), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n1020) );
  XNOR2_X1 U981 ( .A(G160), .B(n1020), .ZN(n908) );
  NAND2_X1 U982 ( .A1(G130), .A2(n885), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G118), .A2(n886), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U985 ( .A1(n889), .A2(G106), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G142), .A2(n724), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  NOR2_X1 U989 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n895), .B(KEYINPUT116), .ZN(n899) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n897) );
  XNOR2_X1 U992 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n903) );
  XNOR2_X1 U995 ( .A(G164), .B(n900), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(n1014), .ZN(n902) );
  XOR2_X1 U997 ( .A(n903), .B(n902), .Z(n906) );
  XOR2_X1 U998 ( .A(n904), .B(G162), .Z(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1001 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT119), .B(n912), .Z(n914) );
  XNOR2_X1 U1004 ( .A(G171), .B(n949), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1006 ( .A(n915), .B(G286), .Z(n916) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n916), .ZN(G397) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2427), .ZN(n926) );
  XOR2_X1 U1009 ( .A(G2430), .B(G2443), .Z(n918) );
  XNOR2_X1 U1010 ( .A(G2435), .B(G2438), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n922) );
  XOR2_X1 U1012 ( .A(G2454), .B(KEYINPUT109), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1015 ( .A(n922), .B(n921), .Z(n924) );
  XNOR2_X1 U1016 ( .A(G2446), .B(KEYINPUT110), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1018 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(n927), .A2(G14), .ZN(n933) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n933), .ZN(n930) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  INV_X1 U1028 ( .A(G96), .ZN(G221) );
  INV_X1 U1029 ( .A(n933), .ZN(G401) );
  XOR2_X1 U1030 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1038) );
  XOR2_X1 U1031 ( .A(KEYINPUT56), .B(G16), .Z(n958) );
  XOR2_X1 U1032 ( .A(G168), .B(G1966), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1034 ( .A(KEYINPUT57), .B(n936), .Z(n948) );
  XNOR2_X1 U1035 ( .A(n937), .B(G1956), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G171), .B(G1961), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G166), .B(G1971), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n940), .B(KEYINPUT123), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n956) );
  XOR2_X1 U1044 ( .A(G1348), .B(n949), .Z(n952) );
  XNOR2_X1 U1045 ( .A(n950), .B(G1341), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n1007) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G22), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G23), .B(G1976), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1055 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n963) );
  XNOR2_X1 U1056 ( .A(n964), .B(n963), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G21), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G5), .B(G1961), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n979) );
  XNOR2_X1 U1061 ( .A(G20), .B(n969), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .Z(n974) );
  XNOR2_X1 U1067 ( .A(G4), .B(n974), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT60), .B(n977), .Z(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1071 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1072 ( .A1(G16), .A2(n981), .ZN(n1004) );
  XOR2_X1 U1073 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1032) );
  XOR2_X1 U1074 ( .A(n1032), .B(KEYINPUT122), .Z(n1001) );
  XNOR2_X1 U1075 ( .A(G2090), .B(G35), .ZN(n996) );
  XOR2_X1 U1076 ( .A(G25), .B(G1991), .Z(n982) );
  NAND2_X1 U1077 ( .A1(n982), .A2(G28), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(G2072), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(G33), .ZN(n991) );
  XOR2_X1 U1080 ( .A(G2067), .B(G26), .Z(n986) );
  INV_X1 U1081 ( .A(G1996), .ZN(n984) );
  XNOR2_X1 U1082 ( .A(n984), .B(G32), .ZN(n985) );
  NAND2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1084 ( .A(G27), .B(n987), .Z(n988) );
  NOR2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(KEYINPUT53), .B(n994), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1090 ( .A(G2084), .B(G34), .Z(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT54), .B(n997), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1001), .B(n1000), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(G29), .A2(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(G11), .A2(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT125), .B(n1008), .Z(n1036) );
  INV_X1 U1099 ( .A(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  XOR2_X1 U1101 ( .A(G160), .B(G2084), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1030) );
  XOR2_X1 U1106 ( .A(G2072), .B(n1020), .Z(n1022) );
  XOR2_X1 U1107 ( .A(G164), .B(G2078), .Z(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT50), .B(n1023), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(G2090), .B(G162), .Z(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT51), .B(n1026), .Z(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(G29), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1119 ( .A(n1038), .B(n1037), .ZN(n1039) );
  XNOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1039), .ZN(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

