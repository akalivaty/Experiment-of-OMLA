//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G250), .B1(G257), .B2(G264), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n207), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n215), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G87), .A2(G250), .ZN(new_n232));
  NAND4_X1  g0032(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n210), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n225), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n202), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n206), .A2(G20), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n217), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n207), .A2(new_n258), .A3(KEYINPUT68), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT68), .B1(new_n207), .B2(new_n258), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G150), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT8), .A2(G58), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT8), .A2(G58), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n258), .A2(G20), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n265), .A2(new_n266), .B1(new_n203), .B2(G20), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n256), .A2(new_n217), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n254), .B1(new_n202), .B2(new_n257), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT9), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n282), .B1(new_n283), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n275), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G190), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n272), .B(new_n289), .C1(new_n290), .C2(new_n288), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n271), .B1(new_n288), .B2(G169), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n259), .A2(new_n260), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n202), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n266), .A2(G77), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n207), .B2(G68), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n269), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n301), .B1(new_n227), .B2(new_n257), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n273), .ZN(new_n311));
  INV_X1    g0111(.A(new_n277), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(G238), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(new_n275), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT13), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(new_n319), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(KEYINPUT14), .B1(new_n321), .B2(G179), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n310), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(G190), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(G200), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n310), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n257), .A2(new_n265), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n252), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT74), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n334), .A3(new_n332), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G58), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n227), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n345), .B2(new_n201), .ZN(new_n346));
  INV_X1    g0146(.A(G159), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n302), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n258), .A3(KEYINPUT3), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT3), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT70), .B1(new_n351), .B2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n207), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n227), .B1(new_n355), .B2(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(KEYINPUT70), .ZN(new_n359));
  AOI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n350), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n348), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n270), .B1(new_n363), .B2(KEYINPUT16), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(new_n348), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n280), .B2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n351), .A2(G33), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n207), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n227), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n366), .B1(new_n373), .B2(KEYINPUT72), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n375), .B(new_n227), .C1(new_n368), .C2(new_n372), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n365), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n343), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n273), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(KEYINPUT75), .A3(new_n273), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G223), .A2(G1698), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n278), .B2(G1698), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n359), .A2(new_n350), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n275), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT76), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n278), .A2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G223), .B2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n354), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n287), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n382), .A4(new_n383), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n290), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n384), .A2(new_n389), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n378), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT17), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n390), .A2(new_n404), .A3(new_n396), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n294), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n343), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n368), .A2(new_n372), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n348), .B1(new_n411), .B2(new_n375), .ZN(new_n412));
  INV_X1    g0212(.A(new_n376), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT16), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n360), .B2(new_n361), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n416));
  OAI211_X1 g0216(.A(KEYINPUT16), .B(new_n366), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n269), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n409), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n408), .A2(new_n419), .A3(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n378), .B2(new_n407), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n403), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g0224(.A(KEYINPUT15), .B(G87), .Z(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n302), .B2(new_n333), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n269), .B1(new_n283), .B2(new_n253), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n257), .A2(new_n283), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n432), .B1(new_n433), .B2(new_n280), .C1(new_n284), .C2(new_n226), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n287), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n311), .B1(new_n312), .B2(G244), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n399), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n431), .B(new_n438), .C1(G200), .C2(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n431), .B1(new_n440), .B2(G169), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n437), .A2(G179), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n298), .A2(new_n330), .A3(new_n424), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT21), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n252), .A2(G116), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT78), .B1(new_n258), .B2(G1), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n206), .A3(G33), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n451), .A3(new_n252), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n269), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n448), .B1(new_n453), .B2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n207), .C1(G33), .C2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n269), .C1(new_n207), .C2(G116), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(KEYINPUT83), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n459), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  INV_X1    g0265(.A(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n206), .B(G45), .C1(new_n466), .C2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT80), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(new_n468), .B1(KEYINPUT5), .B2(new_n466), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(KEYINPUT80), .C1(KEYINPUT5), .C2(new_n466), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n275), .ZN(new_n474));
  INV_X1    g0274(.A(G270), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n465), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(G274), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n287), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G264), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G1698), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G257), .B2(G1698), .ZN(new_n482));
  INV_X1    g0282(.A(G303), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n354), .A2(new_n482), .B1(new_n483), .B2(new_n280), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n477), .A2(new_n479), .B1(new_n484), .B2(new_n287), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n287), .B1(new_n469), .B2(new_n472), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT82), .A3(G270), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n476), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n464), .A2(new_n488), .A3(G169), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n294), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n447), .A2(new_n489), .B1(new_n490), .B2(new_n464), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n488), .A2(G169), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT21), .A4(new_n464), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT84), .B1(new_n489), .B2(new_n447), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n474), .A2(new_n480), .ZN(new_n497));
  INV_X1    g0297(.A(new_n354), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G250), .A3(new_n281), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G257), .A2(G1698), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT88), .B1(new_n354), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  INV_X1    g0303(.A(new_n501), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n359), .A2(new_n503), .A3(new_n350), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n499), .A2(new_n500), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n497), .B1(new_n287), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n477), .A2(new_n479), .ZN(new_n508));
  AOI21_X1  g0308(.A(G169), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n287), .ZN(new_n510));
  INV_X1    g0310(.A(new_n497), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n294), .A2(new_n510), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT89), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n357), .B(new_n369), .C1(KEYINPUT86), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n359), .A2(new_n516), .A3(G87), .A4(new_n350), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  AOI21_X1  g0318(.A(G20), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G87), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n520), .A2(KEYINPUT86), .A3(G20), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n521), .B2(new_n370), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n207), .A2(G107), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT23), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT24), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT87), .B(KEYINPUT24), .C1(new_n519), .C2(new_n525), .ZN(new_n529));
  OR3_X1    g0329(.A1(new_n519), .A2(KEYINPUT24), .A3(new_n525), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n531), .A2(new_n269), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT25), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n252), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n433), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n453), .A2(G107), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n513), .B(new_n514), .C1(new_n532), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n531), .B2(new_n269), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n507), .A2(new_n294), .A3(new_n508), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n510), .A2(new_n511), .A3(new_n508), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G169), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT89), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n496), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n488), .A2(new_n399), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n464), .B1(G200), .B2(new_n488), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(KEYINPUT85), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(KEYINPUT85), .B2(new_n546), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n252), .A2(new_n456), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n453), .B2(new_n456), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(KEYINPUT79), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n410), .A2(G107), .ZN(new_n554));
  XNOR2_X1  g0354(.A(G97), .B(G107), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n558), .A2(G20), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n261), .A2(G77), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n269), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n486), .A2(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n508), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n359), .A2(G244), .A3(new_n350), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(G1698), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n572), .A2(new_n455), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n275), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n576), .A3(new_n294), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n404), .B1(new_n567), .B2(new_n575), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n565), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n568), .A2(new_n576), .A3(G190), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n551), .A2(new_n552), .B1(new_n563), .B2(new_n269), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n567), .B2(new_n575), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n266), .A2(G97), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n207), .B1(new_n316), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n520), .A2(new_n456), .A3(new_n433), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n207), .A2(G68), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n354), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n269), .ZN(new_n592));
  INV_X1    g0392(.A(new_n425), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n253), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n452), .A2(new_n520), .A3(new_n269), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT81), .ZN(new_n597));
  INV_X1    g0397(.A(new_n471), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G250), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n599), .A2(new_n287), .B1(new_n478), .B2(new_n598), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n359), .A2(G238), .A3(new_n281), .A4(new_n350), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n518), .C1(new_n570), .C2(new_n281), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n600), .B1(new_n602), .B2(new_n287), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n595), .B(new_n597), .C1(new_n603), .C2(new_n290), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(G190), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n453), .A2(new_n425), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n592), .A2(new_n606), .A3(new_n594), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n603), .B2(G169), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n603), .A2(new_n294), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n604), .A2(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n584), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n541), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n539), .B(new_n613), .C1(new_n399), .C2(new_n612), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n446), .A2(new_n544), .A3(new_n548), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n609), .ZN(new_n618));
  INV_X1    g0418(.A(new_n608), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  OR3_X1    g0422(.A1(new_n610), .A2(new_n622), .A3(new_n579), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n610), .B2(new_n579), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n539), .A2(new_n542), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n611), .B(new_n614), .C1(new_n496), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n446), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n403), .B(new_n327), .C1(new_n324), .C2(new_n443), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT18), .B1(new_n408), .B2(new_n419), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n378), .A2(new_n407), .A3(new_n421), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT90), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n296), .B1(new_n637), .B2(new_n292), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n629), .A2(new_n638), .ZN(G369));
  NAND3_X1  g0439(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT91), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT91), .ZN(new_n643));
  INV_X1    g0443(.A(G213), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n640), .B2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n464), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n496), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n548), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(KEYINPUT92), .B(G330), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n538), .A2(new_n543), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n614), .ZN(new_n657));
  INV_X1    g0457(.A(new_n648), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n539), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n626), .A2(new_n648), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n496), .A2(new_n658), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n626), .A2(new_n658), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT93), .ZN(G399));
  NOR2_X1   g0470(.A1(new_n212), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n588), .A2(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n221), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  AOI211_X1 g0476(.A(KEYINPUT29), .B(new_n648), .C1(new_n625), .C2(new_n627), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n656), .A2(new_n651), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT96), .A3(new_n616), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT95), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(new_n622), .C1(new_n610), .C2(new_n579), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n621), .B1(new_n683), .B2(new_n623), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT96), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n544), .B2(new_n615), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n679), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n658), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n677), .B1(new_n688), .B2(KEYINPUT29), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n507), .A2(new_n576), .A3(new_n568), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n490), .A4(new_n603), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  INV_X1    g0492(.A(new_n490), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n507), .A2(new_n576), .A3(new_n568), .A4(new_n603), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n603), .B1(new_n568), .B2(new_n576), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n612), .A2(new_n696), .A3(new_n294), .A4(new_n488), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT31), .B1(new_n698), .B2(new_n648), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT94), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n701), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n699), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n616), .A2(new_n544), .A3(new_n548), .A4(new_n658), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n654), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n689), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n676), .B1(new_n709), .B2(G1), .ZN(G364));
  NAND2_X1  g0510(.A1(new_n207), .A2(G13), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n206), .B1(new_n712), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n671), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n212), .A2(new_n370), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G355), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(G116), .B2(new_n211), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n212), .A2(new_n498), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n470), .B2(new_n222), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n247), .A2(new_n470), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(KEYINPUT97), .A2(G169), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n217), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n715), .B1(new_n723), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n290), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n370), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n207), .A2(new_n399), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n294), .A2(new_n290), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G326), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n735), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n483), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n207), .B1(new_n745), .B2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n738), .B(new_n744), .C1(G294), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n294), .A2(G200), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n734), .A2(new_n749), .A3(KEYINPUT98), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT98), .B1(new_n734), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G311), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n734), .A2(new_n745), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G329), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(new_n734), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT33), .B(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n739), .A2(new_n749), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n759), .A2(new_n760), .B1(new_n762), .B2(G322), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n748), .A2(new_n754), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n736), .A2(new_n433), .ZN(new_n765));
  INV_X1    g0565(.A(new_n741), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(G50), .B2(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n767), .B1(new_n344), .B2(new_n761), .C1(new_n752), .C2(new_n283), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n755), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n769));
  INV_X1    g0569(.A(new_n743), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n755), .B2(new_n347), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(new_n280), .A3(new_n772), .ZN(new_n773));
  OR3_X1    g0573(.A1(new_n768), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n758), .A2(new_n227), .B1(new_n746), .B2(new_n456), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n764), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT100), .ZN(new_n778));
  INV_X1    g0578(.A(new_n727), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n777), .B2(KEYINPUT100), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n733), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n730), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n653), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n715), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n655), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n653), .A2(new_n654), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(G396));
  AOI21_X1  g0587(.A(new_n648), .B1(new_n625), .B2(new_n627), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n431), .A2(new_n648), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n439), .A2(new_n790), .B1(new_n442), .B2(new_n441), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n443), .A2(new_n658), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n708), .B(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT105), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n788), .B2(new_n794), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n715), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n798), .B2(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n779), .A2(new_n729), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT101), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n784), .B1(new_n283), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n736), .A2(new_n520), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n743), .A2(new_n433), .B1(new_n755), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n805), .B(new_n807), .C1(G283), .C2(new_n759), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n280), .B1(new_n766), .B2(G303), .ZN(new_n809));
  INV_X1    g0609(.A(G116), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n752), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n761), .A2(new_n812), .B1(new_n746), .B2(new_n456), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT102), .Z(new_n814));
  NOR2_X1   g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  INV_X1    g0616(.A(G150), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n741), .A2(new_n816), .B1(new_n758), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT103), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT104), .B(G143), .Z(new_n820));
  AOI22_X1  g0620(.A1(new_n753), .A2(G159), .B1(new_n762), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(KEYINPUT34), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n736), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G68), .A2(new_n823), .B1(new_n756), .B2(G132), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n202), .B2(new_n743), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n498), .B1(new_n344), .B2(new_n746), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n819), .A2(new_n821), .A3(KEYINPUT34), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n815), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n804), .B1(new_n779), .B2(new_n829), .C1(new_n794), .C2(new_n729), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n800), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NAND3_X1  g0632(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT35), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(G116), .A3(new_n219), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  OR3_X1    g0638(.A1(new_n221), .A2(new_n283), .A3(new_n345), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n202), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n206), .B(G13), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT40), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT108), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n700), .A2(new_n701), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n793), .B1(new_n845), .B2(new_n706), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n648), .B1(new_n309), .B2(new_n308), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n329), .A2(new_n847), .B1(new_n324), .B2(new_n648), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n844), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n846), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n848), .ZN(new_n852));
  NAND2_X1  g0652(.A1(KEYINPUT108), .A2(KEYINPUT40), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  INV_X1    g0655(.A(new_n646), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n419), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n636), .B2(new_n403), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n402), .A3(KEYINPUT90), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n408), .A2(new_n419), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n857), .A3(new_n402), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n857), .A2(new_n402), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n864), .A2(new_n631), .A3(KEYINPUT37), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n855), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n364), .B1(KEYINPUT16), .B2(new_n363), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n336), .B2(new_n335), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n856), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n403), .B2(new_n423), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n408), .B2(new_n856), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .A3(new_n402), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n873), .A2(new_n878), .A3(new_n855), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT106), .B(new_n855), .C1(new_n858), .C2(new_n866), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n869), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n843), .B1(new_n854), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n855), .B1(new_n873), .B2(new_n878), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n846), .A2(new_n849), .A3(new_n853), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT109), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n845), .A2(new_n706), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n446), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n654), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n869), .A2(new_n897), .A3(new_n880), .A4(new_n881), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n324), .A2(new_n658), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT107), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n636), .A2(new_n856), .ZN(new_n905));
  INV_X1    g0705(.A(new_n792), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n788), .B2(new_n794), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(new_n848), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n908), .B2(new_n885), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n901), .B1(new_n898), .B2(new_n899), .ZN(new_n911));
  INV_X1    g0711(.A(new_n907), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n849), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n913), .A2(new_n886), .B1(new_n636), .B2(new_n856), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT107), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n896), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n446), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n689), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n638), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n206), .B2(new_n712), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n917), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n842), .B1(new_n923), .B2(new_n924), .ZN(G367));
  INV_X1    g0725(.A(new_n709), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT114), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n659), .A2(new_n660), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n665), .B1(new_n928), .B2(new_n664), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n661), .B1(new_n655), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n709), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT113), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT113), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n709), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT44), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n579), .A2(new_n658), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n579), .B(new_n583), .C1(new_n581), .C2(new_n658), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n668), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n938), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n665), .A2(new_n666), .A3(new_n939), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n942), .A2(new_n945), .A3(new_n662), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n662), .B1(new_n942), .B2(new_n945), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n927), .B1(new_n935), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n932), .A3(KEYINPUT114), .A4(new_n934), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n926), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n671), .B(KEYINPUT41), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n713), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n595), .A2(new_n597), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n621), .A2(new_n956), .A3(new_n648), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT110), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n610), .B1(new_n956), .B2(new_n648), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT111), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n961), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n657), .A2(new_n664), .A3(new_n939), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n579), .B1(new_n656), .B2(new_n938), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n658), .B2(new_n968), .ZN(new_n969));
  MUX2_X1   g0769(.A(new_n965), .B(new_n963), .S(new_n969), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n661), .A2(new_n939), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n955), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n958), .A2(new_n960), .A3(new_n782), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  NOR4_X1   g0775(.A1(new_n743), .A2(KEYINPUT115), .A3(new_n975), .A4(new_n810), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(KEYINPUT115), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n770), .B2(G116), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(G107), .C2(new_n747), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n753), .A2(G283), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n761), .A2(new_n483), .B1(new_n758), .B2(new_n812), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n741), .A2(new_n806), .B1(new_n755), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n736), .A2(new_n456), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n985), .B(new_n498), .C1(KEYINPUT115), .C2(new_n975), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n979), .A2(new_n980), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n761), .A2(new_n817), .B1(new_n755), .B2(new_n816), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n370), .B(new_n988), .C1(new_n766), .C2(new_n820), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n747), .A2(G68), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n753), .A2(G50), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n736), .A2(new_n283), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n758), .A2(new_n347), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G58), .C2(new_n770), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT47), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n779), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n987), .A2(KEYINPUT47), .A3(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n731), .B1(new_n211), .B2(new_n593), .C1(new_n720), .C2(new_n243), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n715), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n974), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n973), .A2(new_n1003), .ZN(G387));
  OAI211_X1 g0804(.A(new_n935), .B(new_n671), .C1(new_n709), .C2(new_n930), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n930), .A2(new_n714), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n240), .A2(G45), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n673), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n719), .A2(new_n1007), .B1(new_n716), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1010));
  AND3_X1   g0810(.A1(new_n1010), .A2(new_n202), .A3(new_n265), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n673), .B(new_n470), .C1(new_n227), .C2(new_n283), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1010), .B1(new_n202), .B2(new_n265), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1009), .A2(new_n1014), .B1(G107), .B2(new_n211), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n784), .B1(new_n1015), .B2(new_n731), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n593), .A2(new_n746), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n985), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n770), .A2(G77), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1018), .A2(new_n498), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n752), .A2(new_n227), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT117), .B(G150), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1024), .A2(new_n755), .B1(new_n761), .B2(new_n202), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n741), .A2(new_n347), .B1(new_n758), .B2(new_n333), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n752), .A2(new_n483), .B1(new_n982), .B2(new_n761), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT118), .Z(new_n1029));
  INV_X1    g0829(.A(G322), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n806), .B2(new_n758), .C1(new_n1030), .C2(new_n741), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT48), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n770), .A2(G294), .B1(new_n747), .B2(G283), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n736), .A2(new_n810), .B1(new_n755), .B2(new_n742), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n498), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1027), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1016), .B1(new_n928), .B2(new_n782), .C1(new_n1039), .C2(new_n779), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1005), .A2(new_n1006), .A3(new_n1040), .ZN(G393));
  OAI221_X1 g0841(.A(new_n731), .B1(new_n456), .B2(new_n211), .C1(new_n720), .C2(new_n250), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n715), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n202), .A2(new_n758), .B1(new_n743), .B2(new_n227), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n805), .B(new_n1044), .C1(new_n756), .C2(new_n820), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n741), .A2(new_n817), .B1(new_n761), .B2(new_n347), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n753), .A2(new_n265), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n354), .B1(G77), .B2(new_n747), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n741), .A2(new_n982), .B1(new_n761), .B2(new_n806), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT119), .Z(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n280), .B(new_n765), .C1(G116), .C2(new_n747), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n758), .A2(new_n483), .B1(new_n755), .B2(new_n1030), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G283), .B2(new_n770), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n812), .C2(new_n752), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1050), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1043), .B1(new_n1058), .B2(new_n727), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n939), .B2(new_n782), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n948), .B2(new_n713), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n949), .A2(new_n951), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n672), .B1(new_n935), .B2(new_n948), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  NAND3_X1  g0865(.A1(new_n687), .A2(new_n658), .A3(new_n791), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1066), .A2(new_n792), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n901), .B(new_n882), .C1(new_n1067), .C2(new_n848), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n898), .B(new_n899), .C1(new_n902), .C2(new_n908), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n846), .A2(new_n849), .A3(G330), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n707), .A2(new_n849), .A3(new_n654), .A4(new_n794), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1068), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n446), .A2(G330), .A3(new_n891), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n638), .B(new_n1077), .C1(new_n689), .C2(new_n918), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n707), .A2(new_n654), .A3(new_n794), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(new_n848), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n912), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  INV_X1    g0881(.A(G330), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n848), .B1(new_n851), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1067), .A2(new_n1074), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1078), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1086), .A2(KEYINPUT120), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(KEYINPUT120), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1076), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1073), .A2(new_n1075), .A3(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n671), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1076), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n898), .A2(new_n728), .A3(new_n899), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1024), .A2(new_n743), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(KEYINPUT53), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n370), .B(new_n1096), .C1(G50), .C2(new_n823), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1095), .A2(KEYINPUT53), .B1(new_n747), .B2(G159), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  NAND2_X1  g0899(.A1(new_n753), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n758), .A2(new_n816), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G132), .B2(new_n762), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n766), .A2(G128), .B1(new_n756), .B2(G125), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .A4(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G116), .A2(new_n762), .B1(new_n823), .B2(G68), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1106), .A2(new_n370), .A3(new_n771), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n747), .A2(G77), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n753), .A2(G97), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n741), .A2(new_n737), .B1(new_n755), .B2(new_n812), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G107), .B2(new_n759), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n779), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n784), .B(new_n1113), .C1(new_n333), .C2(new_n803), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1092), .A2(new_n714), .B1(new_n1093), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1091), .A2(new_n1115), .ZN(G378));
  NAND2_X1  g0916(.A1(new_n271), .A2(new_n856), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n298), .B(new_n1117), .Z(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1118), .B(new_n1119), .Z(new_n1120));
  AND3_X1   g0920(.A1(new_n910), .A2(new_n915), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n910), .B2(new_n915), .ZN(new_n1122));
  OAI21_X1  g0922(.A(G330), .B1(new_n883), .B2(new_n888), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n887), .B1(new_n852), .B2(new_n844), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n882), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT40), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n888), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1082), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1120), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n904), .B1(new_n903), .B2(new_n909), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT107), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n910), .A2(new_n915), .A3(new_n1120), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n714), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n784), .B1(new_n202), .B2(new_n803), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n466), .B(new_n354), .C1(new_n752), .C2(new_n593), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1020), .B(new_n990), .C1(new_n456), .C2(new_n758), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n741), .A2(new_n810), .B1(new_n761), .B2(new_n433), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n736), .A2(new_n344), .B1(new_n755), .B2(new_n737), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT58), .Z(new_n1144));
  AOI21_X1  g0944(.A(G50), .B1(new_n258), .B2(new_n466), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n498), .B2(G41), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G125), .A2(new_n766), .B1(new_n759), .B2(G132), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n770), .A2(new_n1099), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n762), .A2(G128), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n816), .B2(new_n752), .C1(new_n817), .C2(new_n746), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G33), .B(G41), .C1(new_n756), .C2(G124), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n347), .B2(new_n736), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1144), .B(new_n1146), .C1(new_n1152), .C2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n727), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1138), .B1(new_n1159), .B2(new_n1161), .C1(new_n1120), .C2(new_n729), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT123), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1137), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1123), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1078), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1090), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1133), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .A4(KEYINPUT57), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n672), .B1(new_n1173), .B2(KEYINPUT124), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT124), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1136), .A2(new_n1175), .A3(KEYINPUT57), .A4(new_n1167), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT125), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1172), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1176), .A3(KEYINPUT125), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1164), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G375));
  NAND3_X1  g0982(.A1(new_n1081), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n953), .B(new_n1183), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n761), .A2(new_n737), .B1(new_n758), .B2(new_n810), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1017), .A2(new_n1185), .A3(new_n280), .A4(new_n992), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G97), .A2(new_n770), .B1(new_n756), .B2(G303), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n812), .B2(new_n741), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G107), .B2(new_n753), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G132), .A2(new_n766), .B1(new_n762), .B2(G137), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n759), .A2(new_n1099), .B1(new_n756), .B2(G128), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G150), .B2(new_n753), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n743), .A2(new_n347), .B1(new_n736), .B2(new_n344), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n354), .B(new_n1194), .C1(G50), .C2(new_n747), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1186), .A2(new_n1189), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n715), .B1(G68), .B2(new_n802), .C1(new_n1196), .C2(new_n779), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n848), .B2(new_n728), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n714), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1184), .A2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(G378), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1181), .A2(new_n1202), .ZN(new_n1203));
  OR4_X1    g1003(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1204));
  OR4_X1    g1004(.A1(G387), .A2(new_n1203), .A3(G390), .A4(new_n1204), .ZN(G407));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1203), .ZN(G409));
  NAND2_X1  g1006(.A1(G387), .A2(new_n1064), .ZN(new_n1207));
  XOR2_X1   g1007(.A(G393), .B(G396), .Z(new_n1208));
  NAND3_X1  g1008(.A1(new_n973), .A2(new_n1003), .A3(G390), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1208), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G390), .B1(new_n973), .B2(new_n1003), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1002), .B(new_n1064), .C1(new_n955), .C2(new_n972), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  AND4_X1   g1015(.A1(new_n1091), .A2(new_n1137), .A3(new_n1115), .A4(new_n1162), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1136), .A2(new_n953), .A3(new_n1167), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1216), .A2(new_n1217), .B1(G213), .B2(new_n647), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1181), .B2(new_n1202), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT60), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n672), .B(new_n1085), .C1(new_n1220), .C2(new_n1183), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1220), .B2(new_n1183), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1222), .A2(G384), .A3(new_n1200), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G384), .B1(new_n1222), .B2(new_n1200), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n647), .A2(G213), .A3(G2897), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT126), .Z(new_n1227));
  XNOR2_X1  g1027(.A(new_n1225), .B(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(KEYINPUT61), .B(new_n1215), .C1(new_n1219), .C2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1218), .B(new_n1225), .C1(new_n1181), .C2(new_n1202), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT127), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1180), .A3(new_n1171), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1164), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1202), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1218), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(KEYINPUT63), .A4(new_n1225), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1230), .A2(KEYINPUT62), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1174), .A2(new_n1176), .A3(KEYINPUT125), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT125), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1172), .ZN(new_n1246));
  OAI21_X1  g1046(.A(G378), .B1(new_n1246), .B2(new_n1164), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1218), .A4(new_n1225), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1228), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1243), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1215), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1242), .A2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1203), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1225), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1215), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1247), .B(new_n1203), .C1(new_n1224), .C2(new_n1223), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(G402));
endmodule


