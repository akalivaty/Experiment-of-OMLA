//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT75), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n207), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n213), .ZN(new_n216));
  AND2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT76), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT76), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n220), .A3(new_n206), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n214), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT69), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(G120gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n227), .B2(G120gat), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n237));
  INV_X1    g036(.A(G134gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G127gat), .ZN(new_n239));
  INV_X1    g038(.A(G127gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G134gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n237), .A2(new_n239), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n227), .A2(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n239), .A2(new_n241), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n239), .B2(new_n241), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n224), .A2(new_n226), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n241), .A3(new_n251), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n258), .A2(new_n259), .B1(new_n249), .B2(new_n248), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n233), .A2(new_n235), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n243), .B1(new_n261), .B2(new_n231), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n214), .A2(new_n222), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n245), .A2(new_n254), .A3(new_n214), .A4(new_n222), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G225gat), .A2(G233gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n256), .A2(new_n265), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n223), .B1(new_n260), .B2(new_n262), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  INV_X1    g072(.A(new_n269), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n267), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n264), .A2(new_n254), .A3(new_n245), .A4(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n277), .A2(new_n279), .A3(new_n271), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n223), .A2(KEYINPUT3), .B1(new_n245), .B2(new_n254), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n281), .B2(new_n226), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n270), .A2(new_n275), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT80), .ZN(new_n285));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n287), .B(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n275), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n282), .A2(new_n271), .A3(new_n279), .A4(new_n277), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n290), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(KEYINPUT6), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT83), .B(G22gat), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(G211gat), .A2(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307));
  AND2_X1   g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n304), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n314), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n223), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n303), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n226), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n315), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n324), .B(new_n317), .C1(new_n318), .C2(new_n303), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n302), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT31), .B(G50gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n326), .A2(G22gat), .A3(new_n327), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n326), .A2(new_n327), .A3(new_n302), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n328), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT84), .B(new_n302), .C1(new_n326), .C2(new_n327), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n332), .B(KEYINPUT81), .Z(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT64), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(KEYINPUT64), .A3(new_n345), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT23), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT25), .A2(new_n357), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n346), .A2(new_n351), .A3(new_n352), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT27), .B(G183gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n350), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n349), .A2(KEYINPUT27), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G183gat), .ZN(new_n373));
  AND4_X1   g172(.A1(new_n368), .A2(new_n371), .A3(new_n373), .A4(new_n350), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT65), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT65), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n355), .A3(new_n356), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n377), .A2(new_n360), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n344), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n382), .B2(new_n344), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n367), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT72), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n320), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(new_n344), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT66), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n384), .A3(new_n375), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n367), .A3(new_n389), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n391), .A2(new_n322), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n322), .B1(new_n391), .B2(new_n395), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n343), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n395), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n394), .A2(new_n367), .B1(new_n320), .B2(new_n389), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n323), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n391), .A2(new_n322), .A3(new_n395), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT73), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT74), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n398), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT30), .A4(new_n407), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n401), .A2(new_n402), .A3(new_n407), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT40), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n256), .A2(new_n277), .A3(new_n279), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT39), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n274), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n290), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n272), .A2(new_n266), .A3(new_n269), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT39), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n274), .B2(new_n416), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n274), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT39), .A3(new_n420), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(KEYINPUT40), .A3(new_n290), .A4(new_n418), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n290), .B1(new_n294), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n428), .B2(new_n294), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n295), .B1(new_n283), .B2(KEYINPUT85), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n294), .A2(new_n428), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n291), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT37), .B1(new_n396), .B2(new_n397), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n402), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n408), .A4(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n434), .A2(new_n298), .A3(new_n411), .A4(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n437), .A2(new_n408), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n398), .A2(new_n403), .A3(KEYINPUT37), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n342), .B(new_n431), .C1(new_n440), .C2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n413), .A2(new_n410), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n299), .A2(new_n445), .A3(new_n409), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n337), .A2(new_n336), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n329), .ZN(new_n448));
  INV_X1    g247(.A(new_n339), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n341), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n335), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n387), .A2(new_n263), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n367), .B(new_n255), .C1(new_n385), .C2(new_n386), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G15gat), .B(G43gat), .Z(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n458), .B(KEYINPUT32), .C1(new_n460), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n454), .A2(new_n457), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n455), .ZN(new_n470));
  AOI211_X1 g269(.A(KEYINPUT34), .B(new_n456), .C1(new_n454), .C2(new_n457), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n457), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n255), .B1(new_n394), .B2(new_n367), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n455), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT34), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n468), .A3(new_n455), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT71), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n465), .B(new_n467), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n467), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(KEYINPUT71), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n444), .A2(new_n453), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n480), .B(new_n483), .C1(new_n450), .C2(new_n451), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT35), .B1(new_n489), .B2(new_n446), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n409), .A2(new_n491), .A3(new_n410), .A4(new_n413), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n298), .B2(new_n434), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n480), .A2(new_n483), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n342), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n488), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G8gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT90), .B(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n513), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(KEYINPUT15), .A3(new_n514), .A4(new_n515), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n510), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n510), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n528), .A4(new_n530), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n510), .B(new_n523), .Z(new_n535));
  XOR2_X1   g334(.A(new_n528), .B(KEYINPUT13), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT89), .B(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT11), .B(G169gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT12), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n533), .A2(new_n534), .A3(new_n537), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n531), .A2(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(KEYINPUT92), .A3(new_n534), .A4(new_n543), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n534), .ZN(new_n550));
  INV_X1    g349(.A(new_n543), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n498), .A2(new_n500), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT93), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n498), .A2(new_n556), .A3(new_n500), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559));
  XOR2_X1   g358(.A(G57gat), .B(G64gat), .Z(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  NAND3_X1  g372(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n577), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n559), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT101), .Z(new_n581));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(new_n587), .A3(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n578), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n579), .B2(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT100), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n579), .A2(new_n587), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n578), .A4(new_n588), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n559), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n559), .B(KEYINPUT102), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n594), .A2(new_n578), .A3(new_n600), .A4(new_n588), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT103), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n588), .A2(new_n578), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(KEYINPUT103), .A3(new_n600), .A4(new_n594), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n585), .B1(new_n606), .B2(new_n581), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT104), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n598), .A2(new_n610), .A3(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n577), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n524), .B2(new_n526), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n523), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT97), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT95), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n615), .A2(new_n620), .A3(new_n617), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n623), .A2(new_n624), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n628), .B(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n636));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  AOI21_X1  g437(.A(new_n529), .B1(KEYINPUT21), .B2(new_n567), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT94), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n640), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n613), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT105), .B1(new_n558), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n651), .B(new_n652), .C1(new_n555), .C2(new_n557), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n300), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  OAI211_X1 g455(.A(new_n414), .B(new_n656), .C1(new_n650), .C2(new_n653), .ZN(new_n657));
  INV_X1    g456(.A(new_n414), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n558), .A2(new_n649), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n651), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n558), .A2(KEYINPUT105), .A3(new_n649), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(new_n509), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT42), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n668), .B(new_n494), .C1(new_n650), .C2(new_n653), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n485), .A2(new_n487), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n660), .B2(new_n661), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n669), .B1(new_n674), .B2(new_n668), .ZN(G1326gat));
  OAI21_X1  g474(.A(new_n452), .B1(new_n650), .B2(new_n653), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT107), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n678), .B(new_n452), .C1(new_n650), .C2(new_n653), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n677), .B2(new_n679), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n613), .A2(new_n647), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n635), .B(new_n685), .C1(new_n555), .C2(new_n557), .ZN(new_n686));
  INV_X1    g485(.A(G29gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n300), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n671), .A2(new_n453), .A3(new_n444), .A4(new_n672), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n635), .B1(new_n692), .B2(new_n496), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n498), .A2(KEYINPUT44), .A3(new_n500), .A4(new_n634), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n553), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n685), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n696), .A2(new_n300), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n690), .B(new_n691), .C1(new_n687), .C2(new_n699), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n658), .A2(new_n511), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n686), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n702), .A2(KEYINPUT108), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(new_n414), .A3(new_n698), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n511), .B1(new_n702), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n702), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n673), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n709), .A3(new_n695), .A4(new_n698), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n484), .A2(G43gat), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n710), .A2(G43gat), .B1(new_n686), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1330gat));
  NAND4_X1  g513(.A1(new_n696), .A2(G50gat), .A3(new_n452), .A4(new_n698), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n686), .A2(new_n452), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(G50gat), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT48), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n715), .B(new_n719), .C1(G50gat), .C2(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1331gat));
  NAND2_X1  g520(.A1(new_n692), .A2(new_n496), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n648), .A2(new_n612), .A3(new_n553), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT110), .Z(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n300), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g526(.A(new_n724), .B(KEYINPUT110), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n658), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  NAND3_X1  g532(.A1(new_n725), .A2(new_n562), .A3(new_n494), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n728), .A2(new_n673), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n562), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(KEYINPUT50), .C1(new_n562), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n728), .A2(new_n342), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n563), .ZN(G1335gat));
  NOR3_X1   g541(.A1(new_n612), .A2(new_n553), .A3(new_n647), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n696), .A2(new_n300), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n553), .A2(new_n647), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n693), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n693), .A2(KEYINPUT51), .A3(new_n745), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n746), .A2(KEYINPUT111), .A3(new_n747), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n613), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n300), .A2(new_n569), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n744), .A2(new_n569), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n694), .A2(new_n414), .A3(new_n695), .A4(new_n743), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n658), .A2(G92gat), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n756), .B(new_n758), .C1(new_n753), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n748), .A2(KEYINPUT112), .A3(new_n750), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n763), .A3(new_n747), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n762), .A2(new_n613), .A3(new_n764), .A4(new_n759), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n758), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n766), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n696), .A2(new_n709), .A3(new_n743), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G99gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n752), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n612), .A2(G99gat), .A3(new_n484), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT113), .Z(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n753), .A2(G106gat), .A3(new_n342), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n694), .A2(new_n452), .A3(new_n695), .A4(new_n743), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n612), .A2(G106gat), .A3(new_n342), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n764), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n776), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n774), .A2(new_n778), .B1(new_n781), .B2(new_n777), .ZN(G1339gat));
  INV_X1    g581(.A(new_n647), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n606), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n594), .A2(new_n578), .A3(new_n588), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(new_n599), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n597), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n785), .A2(KEYINPUT55), .A3(new_n585), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n584), .B1(new_n606), .B2(new_n784), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT55), .A4(new_n788), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n785), .A2(new_n585), .A3(new_n788), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n794), .A2(new_n634), .A3(new_n598), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n535), .A2(new_n536), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n542), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n549), .A2(KEYINPUT115), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT115), .B1(new_n549), .B2(new_n801), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n794), .A2(new_n553), .A3(new_n598), .A4(new_n797), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n609), .A2(new_n549), .A3(new_n611), .A4(new_n801), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n634), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n783), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n649), .A2(new_n697), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n299), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n658), .A2(new_n811), .A3(new_n342), .A4(new_n494), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n553), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n228), .B2(new_n230), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n227), .B2(new_n813), .ZN(G1340gat));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n613), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n647), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G127gat), .ZN(G1342gat));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n812), .B(new_n634), .C1(new_n820), .C2(new_n238), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n238), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n807), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n635), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n634), .A2(new_n598), .A3(new_n797), .ZN(new_n827));
  INV_X1    g626(.A(new_n804), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n794), .A4(new_n802), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n647), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n810), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n824), .B(new_n300), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n709), .A2(new_n414), .A3(new_n342), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n811), .A2(new_n824), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n553), .A2(new_n202), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT119), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n299), .A2(new_n414), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n673), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n342), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n795), .A2(KEYINPUT116), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n791), .A2(new_n847), .A3(new_n788), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n796), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(new_n794), .A3(new_n553), .A4(new_n598), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n807), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n635), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n647), .B1(new_n852), .B2(new_n829), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n843), .B(new_n845), .C1(new_n853), .C2(new_n831), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n342), .B1(new_n809), .B2(new_n810), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(KEYINPUT57), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n634), .B1(new_n850), .B2(new_n807), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n783), .B1(new_n857), .B2(new_n805), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n810), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n843), .B1(new_n859), .B2(new_n845), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n553), .B(new_n842), .C1(new_n856), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n839), .B1(new_n861), .B2(G141gat), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n863), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n865), .B(new_n839), .C1(new_n861), .C2(G141gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(G1344gat));
  NOR2_X1   g666(.A1(new_n834), .A2(new_n835), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n203), .A3(new_n613), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G148gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n860), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n841), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n873), .B2(new_n613), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n809), .A2(new_n810), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n452), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n844), .A3(new_n452), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n877), .A2(new_n613), .A3(new_n842), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n870), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n869), .B1(new_n874), .B2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n868), .A2(new_n208), .A3(new_n647), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n872), .A2(new_n783), .A3(new_n841), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n208), .ZN(G1346gat));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n209), .A3(new_n634), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n872), .A2(new_n635), .A3(new_n841), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n209), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n489), .A2(new_n300), .A3(new_n658), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n875), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n355), .A3(new_n697), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(KEYINPUT121), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n553), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n355), .ZN(G1348gat));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n356), .A3(new_n613), .ZN(new_n894));
  OAI21_X1  g693(.A(G176gat), .B1(new_n889), .B2(new_n612), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1349gat));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n647), .A2(new_n369), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n889), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G183gat), .B1(new_n889), .B2(new_n783), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n889), .B2(new_n898), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n903));
  NAND2_X1  g702(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT124), .Z(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n902), .B(new_n905), .C1(KEYINPUT123), .C2(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n889), .B2(new_n635), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT61), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n350), .A3(new_n634), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n300), .A2(new_n658), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n877), .A2(new_n673), .A3(new_n878), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n697), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n855), .A2(new_n673), .A3(new_n914), .ZN(new_n918));
  INV_X1    g717(.A(G197gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n553), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1352gat));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n918), .A2(new_n924), .A3(new_n925), .A4(new_n613), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n915), .B2(new_n612), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n925), .A3(new_n613), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n928), .B(new_n929), .C1(new_n932), .C2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n310), .A3(new_n647), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n915), .A2(new_n783), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT63), .B(G211gat), .C1(new_n915), .C2(new_n783), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n937), .B2(new_n939), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n915), .B2(new_n635), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n918), .A2(new_n311), .A3(new_n634), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1355gat));
endmodule


