//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT64), .B(G238), .Z(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n218), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n220), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n243), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G274), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n251), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(G244), .ZN(new_n260));
  INV_X1    g0060(.A(G179), .ZN(new_n261));
  INV_X1    g0061(.A(new_n251), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G107), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n219), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(G232), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n271), .A2(new_n272), .A3(G1698), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n262), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n260), .A2(new_n261), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n213), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n206), .A2(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G77), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n278), .A2(new_n280), .B1(G77), .B2(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G20), .A2(G77), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G87), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT15), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G87), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n207), .A2(G33), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n282), .B1(new_n283), .B2(new_n285), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n277), .A2(new_n213), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n260), .A2(new_n274), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT71), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n275), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI211_X1 g0100(.A(KEYINPUT71), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT69), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT69), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n260), .A2(new_n306), .A3(new_n274), .A4(G190), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT70), .B(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(new_n295), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(G150), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n283), .A2(new_n292), .B1(new_n313), .B2(new_n285), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G20), .B2(new_n203), .ZN(new_n315));
  INV_X1    g0115(.A(new_n294), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n279), .A2(G50), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n278), .A2(new_n318), .B1(G50), .B2(new_n276), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n269), .A2(G222), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n323), .B2(new_n269), .C1(new_n324), .C2(new_n267), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n262), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT67), .B(G226), .Z(new_n327));
  AOI21_X1  g0127(.A(new_n254), .B1(new_n259), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G179), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n320), .B(new_n330), .C1(new_n297), .C2(new_n329), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n317), .A2(new_n319), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n320), .A2(KEYINPUT9), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n326), .A2(G190), .A3(new_n328), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(new_n308), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n334), .A2(new_n335), .A3(new_n338), .A4(new_n339), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n331), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n303), .A2(new_n344), .A3(new_n310), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n312), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n283), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n279), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n348), .A2(new_n278), .B1(new_n276), .B2(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT78), .ZN(new_n350));
  INV_X1    g0150(.A(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n220), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n284), .A2(G159), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT7), .B1(new_n271), .B2(new_n207), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n357), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT77), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n357), .B1(new_n269), .B2(G20), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n265), .A2(G33), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT7), .B(new_n207), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AOI211_X1 g0165(.A(new_n360), .B(new_n220), .C1(new_n362), .C2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT16), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n355), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n294), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n350), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n220), .B1(new_n362), .B2(new_n365), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n369), .B1(new_n374), .B2(KEYINPUT77), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n371), .B1(new_n375), .B2(new_n366), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n355), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n316), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n349), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n269), .A2(G223), .A3(new_n321), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  INV_X1    g0182(.A(G226), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n267), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n262), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n255), .A2(new_n272), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n254), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n261), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n297), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT18), .B1(new_n380), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n349), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n378), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT78), .B1(new_n376), .B2(new_n378), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n393), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G190), .B2(new_n391), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n395), .B(new_n404), .C1(new_n396), .C2(new_n397), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n373), .A2(new_n379), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n395), .A4(new_n404), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n394), .A2(new_n401), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n254), .B1(new_n259), .B2(G238), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n264), .A2(new_n266), .A3(G232), .A4(G1698), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(new_n321), .ZN(new_n415));
  AND3_X1   g0215(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n262), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n412), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n258), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n257), .B1(new_n251), .B2(new_n253), .ZN(new_n423));
  OAI21_X1  g0223(.A(G238), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n254), .ZN(new_n425));
  AND4_X1   g0225(.A1(new_n412), .A2(new_n424), .A3(new_n420), .A4(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n413), .A2(new_n412), .A3(new_n420), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT74), .ZN(new_n433));
  INV_X1    g0233(.A(new_n421), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n413), .A2(new_n435), .A3(new_n412), .A4(new_n420), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(G179), .A4(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(G169), .B1(new_n428), .B2(new_n429), .C1(new_n421), .C2(new_n426), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n323), .B2(new_n292), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n294), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT11), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT75), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(KEYINPUT75), .A3(new_n445), .ZN(new_n449));
  INV_X1    g0249(.A(new_n276), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n220), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT12), .ZN(new_n452));
  INV_X1    g0252(.A(new_n278), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G68), .A3(new_n279), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n448), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n439), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n433), .A2(new_n434), .A3(G190), .A4(new_n436), .ZN(new_n458));
  INV_X1    g0258(.A(new_n456), .ZN(new_n459));
  OAI21_X1  g0259(.A(G200), .B1(new_n421), .B2(new_n426), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n346), .A2(KEYINPUT80), .A3(new_n411), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(new_n312), .A3(new_n343), .A4(new_n345), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n410), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n264), .A2(new_n266), .A3(G250), .A4(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(new_n321), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n262), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(G274), .A3(new_n251), .A4(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(new_n251), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G257), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n474), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n297), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n470), .A2(new_n471), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .A4(new_n321), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n468), .A4(new_n469), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n488), .A2(new_n262), .B1(G257), .B2(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n261), .A3(new_n478), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n491), .A2(new_n492), .A3(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(G97), .B(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n495), .A2(new_n207), .B1(new_n323), .B2(new_n285), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n268), .B1(new_n362), .B2(new_n365), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n294), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n276), .A2(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n278), .B1(new_n206), .B2(G33), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n485), .A2(new_n490), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n474), .A2(G190), .A3(new_n478), .A4(new_n483), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n498), .A3(new_n501), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n402), .B1(new_n489), .B2(new_n478), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n501), .ZN(new_n509));
  INV_X1    g0309(.A(new_n497), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n494), .A2(new_n491), .ZN(new_n511));
  INV_X1    g0311(.A(new_n493), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n515), .B2(new_n294), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n484), .A2(G200), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT81), .A4(new_n505), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n503), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n264), .A2(new_n266), .A3(new_n207), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n269), .A2(new_n523), .A3(new_n207), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n292), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n207), .B2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n528), .B(new_n531), .C1(new_n207), .C2(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n525), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n316), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n453), .B1(G1), .B2(new_n263), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT25), .B1(new_n450), .B2(new_n268), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n450), .A2(KEYINPUT25), .A3(new_n268), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n539), .A2(new_n268), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n481), .A2(G264), .A3(new_n251), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n478), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n269), .A2(G250), .A3(new_n321), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n262), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n261), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G169), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n520), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n262), .ZN(new_n554));
  INV_X1    g0354(.A(new_n545), .ZN(new_n555));
  AOI21_X1  g0355(.A(G169), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n261), .B2(new_n550), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(KEYINPUT86), .C1(new_n538), .C2(new_n542), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(G190), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n543), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n553), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n500), .A2(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n450), .A2(new_n526), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n277), .A2(new_n213), .B1(G20), .B2(new_n526), .ZN(new_n567));
  AOI21_X1  g0367(.A(G20), .B1(G33), .B2(G283), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n263), .A2(G97), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT84), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT84), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(KEYINPUT20), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n481), .A2(G270), .A3(new_n251), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n478), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n269), .A2(G264), .A3(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n269), .A2(G257), .A3(new_n321), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n271), .A2(G303), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n262), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G190), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n576), .B(new_n584), .C1(new_n402), .C2(new_n583), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n262), .ZN(new_n587));
  INV_X1    g0387(.A(new_n578), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G169), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n586), .B1(new_n576), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n574), .A2(new_n575), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n565), .A3(new_n564), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(G179), .A3(new_n583), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(KEYINPUT21), .A3(G169), .A4(new_n589), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n585), .A2(new_n591), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n267), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n264), .A2(new_n266), .A3(G238), .A4(new_n321), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n269), .A2(new_n601), .A3(G238), .A4(new_n321), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n251), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n477), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n605), .A2(G250), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n251), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n252), .B2(new_n605), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n261), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n269), .A2(new_n207), .A3(G68), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n292), .A2(new_n492), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(KEYINPUT19), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT19), .B1(new_n416), .B2(new_n417), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G97), .A2(G107), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n207), .B1(new_n286), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n294), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n291), .A2(new_n450), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n500), .A2(new_n290), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n618), .A4(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n297), .B1(new_n604), .B2(new_n608), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n610), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n609), .A2(G190), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n500), .A2(G87), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n617), .A2(new_n618), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n308), .B1(new_n604), .B2(new_n608), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n596), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n467), .A2(new_n519), .A3(new_n563), .A4(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n630), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT87), .B(new_n297), .C1(new_n604), .C2(new_n608), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n610), .A2(new_n637), .A3(new_n620), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n519), .A3(new_n562), .ZN(new_n640));
  INV_X1    g0440(.A(new_n543), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n557), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT88), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n639), .A2(new_n646), .A3(new_n503), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n638), .A2(new_n636), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n625), .A2(new_n503), .A3(new_n630), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n467), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n457), .B1(new_n653), .B2(new_n302), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n407), .A2(new_n409), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n394), .B(new_n401), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n340), .A2(new_n342), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n331), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(G369));
  XOR2_X1   g0459(.A(new_n643), .B(KEYINPUT88), .Z(new_n660));
  NAND3_X1  g0460(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n576), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n596), .A2(new_n667), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n668), .A2(KEYINPUT89), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT89), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n563), .B1(new_n543), .B2(new_n665), .ZN(new_n675));
  INV_X1    g0475(.A(new_n642), .ZN(new_n676));
  INV_X1    g0476(.A(new_n665), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n563), .A2(new_n643), .A3(new_n665), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n676), .B2(new_n665), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n615), .A2(new_n286), .A3(new_n526), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n206), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n217), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  OAI21_X1  g0490(.A(new_n665), .B1(new_n645), .B2(new_n651), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n694));
  AOI211_X1 g0494(.A(KEYINPUT92), .B(new_n503), .C1(new_n508), .C2(new_n518), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n508), .A2(new_n518), .ZN(new_n697));
  INV_X1    g0497(.A(new_n503), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n639), .A2(new_n562), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n553), .A2(new_n558), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(new_n643), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n648), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n639), .A2(new_n503), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(KEYINPUT26), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n677), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n691), .A2(new_n710), .A3(new_n692), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n694), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n609), .A2(new_n489), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n550), .A2(new_n583), .A3(G179), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n550), .A2(new_n583), .A3(G179), .ZN(new_n717));
  INV_X1    g0517(.A(new_n609), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n484), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n587), .A2(new_n588), .A3(G179), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n560), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n489), .A4(new_n609), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n723), .B2(new_n677), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n716), .A2(new_n719), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n716), .A2(new_n719), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n563), .A2(new_n632), .A3(new_n519), .A4(new_n665), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n673), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n712), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n690), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n206), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n686), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n674), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n672), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(G330), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n213), .B1(G20), .B2(new_n297), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n207), .A2(new_n261), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n754), .A2(new_n402), .A3(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G68), .B1(G77), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n754), .A2(new_n304), .A3(new_n402), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n754), .A2(new_n304), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n759), .B1(new_n202), .B2(new_n761), .C1(new_n351), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n308), .A2(new_n304), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(G107), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n756), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n207), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n492), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n308), .A2(G190), .A3(new_n765), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n271), .B1(new_n778), .B2(G87), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(KEYINPUT93), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(KEYINPUT93), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n768), .A2(new_n776), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n269), .B(new_n784), .C1(G326), .C2(new_n760), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G311), .A2(new_n758), .B1(new_n770), .B2(G329), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n755), .A2(new_n787), .B1(new_n762), .B2(G322), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n790), .A2(new_n766), .B1(new_n777), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n782), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n752), .B1(new_n793), .B2(KEYINPUT94), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(KEYINPUT94), .B2(new_n793), .ZN(new_n795));
  INV_X1    g0595(.A(new_n742), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n210), .A2(G355), .A3(new_n269), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n685), .A2(new_n269), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n216), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n248), .A2(new_n476), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(G116), .B2(new_n210), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n748), .A2(new_n751), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n745), .B1(new_n750), .B2(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n295), .A2(new_n665), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n310), .B(new_n807), .C1(new_n300), .C2(new_n301), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n298), .A2(new_n299), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n298), .A2(new_n299), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n809), .A2(new_n810), .A3(new_n275), .A4(new_n806), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n691), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n812), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n665), .C1(new_n645), .C2(new_n651), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n742), .B1(new_n816), .B2(new_n734), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n734), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n751), .A2(new_n746), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n742), .B1(new_n820), .B2(G77), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n763), .A2(new_n783), .B1(new_n757), .B2(new_n526), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n761), .A2(new_n791), .B1(new_n769), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n269), .B(new_n775), .C1(G283), .C2(new_n755), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n767), .A2(G87), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n778), .A2(G107), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n762), .A2(G143), .B1(G159), .B2(new_n758), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(new_n755), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n761), .C1(new_n313), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT34), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n767), .A2(G68), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n778), .A2(G50), .ZN(new_n836));
  INV_X1    g0636(.A(new_n774), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G58), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n271), .B1(new_n770), .B2(G132), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n829), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n821), .B1(new_n841), .B2(new_n751), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n814), .B2(new_n747), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n818), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n739), .A2(new_n206), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n398), .A2(new_n399), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n398), .A2(new_n664), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n405), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n395), .B1(new_n372), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n399), .B2(new_n664), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n405), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n850), .B1(new_n854), .B2(new_n849), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n852), .A2(new_n664), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n410), .A2(KEYINPUT96), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT96), .B1(new_n410), .B2(new_n856), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n855), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n847), .A2(new_n848), .A3(new_n405), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n850), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n410), .A2(new_n398), .A3(new_n664), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n860), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n439), .A2(new_n456), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(new_n677), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n863), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n664), .B1(new_n394), .B2(new_n401), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n861), .A2(new_n862), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n456), .A2(new_n677), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(new_n653), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n456), .B(new_n677), .C1(new_n461), .C2(new_n439), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n303), .A2(new_n677), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n815), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n876), .B1(new_n877), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n875), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n694), .A2(new_n467), .A3(new_n711), .A4(new_n709), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n888), .A2(new_n658), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n724), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n732), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n812), .B1(new_n879), .B2(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT98), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n891), .B1(new_n897), .B2(new_n870), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT97), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT97), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n891), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n862), .B2(new_n861), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n467), .A2(new_n894), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n673), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n846), .B1(new_n890), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n890), .B2(new_n907), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n910), .A2(G116), .A3(new_n214), .A4(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OAI21_X1  g0713(.A(G77), .B1(new_n351), .B2(new_n220), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n244), .B1(new_n216), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n738), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(G367));
  INV_X1    g0717(.A(KEYINPUT101), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n639), .B1(new_n628), .B2(new_n665), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n628), .A2(new_n665), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n648), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT43), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n698), .A2(new_n665), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n502), .A2(new_n677), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n700), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT42), .B1(new_n925), .B2(new_n681), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n697), .A2(new_n698), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT92), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n519), .A2(new_n696), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n924), .ZN(new_n930));
  INV_X1    g0730(.A(new_n923), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n933), .A3(new_n682), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT99), .ZN(new_n935));
  INV_X1    g0735(.A(new_n702), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n698), .C1(new_n930), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n665), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n700), .A2(new_n702), .A3(new_n924), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n935), .B1(new_n939), .B2(new_n698), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n926), .B(new_n934), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT100), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n933), .B1(new_n932), .B2(new_n682), .ZN(new_n944));
  AOI211_X1 g0744(.A(KEYINPUT42), .B(new_n681), .C1(new_n930), .C2(new_n931), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n698), .B1(new_n930), .B2(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT99), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n665), .A3(new_n937), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT100), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n918), .B(new_n922), .C1(new_n943), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n942), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT100), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n953), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n918), .B1(new_n957), .B2(new_n922), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT102), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n680), .A2(new_n925), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n962), .A2(KEYINPUT103), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT103), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n962), .A2(new_n963), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT103), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(KEYINPUT103), .A3(new_n963), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n960), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n740), .B(KEYINPUT106), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n683), .A2(new_n932), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  INV_X1    g0774(.A(new_n683), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n925), .C1(KEYINPUT104), .C2(KEYINPUT44), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n683), .C2(new_n932), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n976), .B(new_n979), .C1(new_n977), .C2(new_n978), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n974), .A2(new_n680), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n680), .B1(new_n980), .B2(new_n974), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n681), .A2(KEYINPUT105), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n679), .B1(new_n643), .B2(new_n665), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n681), .A2(KEYINPUT105), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n674), .B(new_n987), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n735), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n686), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n972), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n966), .A2(new_n971), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n798), .A2(new_n239), .ZN(new_n993));
  INV_X1    g0793(.A(new_n802), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n685), .B2(new_n290), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n796), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G283), .A2(new_n758), .B1(new_n770), .B2(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n763), .B2(new_n791), .C1(new_n823), .C2(new_n761), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n777), .A2(new_n526), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n271), .B1(new_n268), .B2(new_n774), .C1(new_n832), .C2(new_n783), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n766), .A2(new_n492), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT107), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n271), .B1(new_n760), .B2(G143), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n220), .B2(new_n774), .ZN(new_n1006));
  INV_X1    g0806(.A(G159), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n313), .A2(new_n763), .B1(new_n832), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n757), .A2(new_n202), .B1(new_n769), .B2(new_n831), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n351), .B2(new_n777), .C1(new_n323), .C2(new_n766), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n996), .B1(new_n749), .B2(new_n921), .C1(new_n1013), .C2(new_n752), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n992), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n972), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n675), .A2(new_n678), .A3(new_n748), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n210), .A2(new_n269), .A3(new_n687), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(G107), .B2(new_n210), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n236), .A2(G45), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n283), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n685), .B(new_n269), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n742), .B1(new_n1025), .B2(new_n994), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT108), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n269), .B1(new_n769), .B2(new_n313), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1028), .B(new_n1002), .C1(G77), .C2(new_n778), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT109), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n774), .A2(new_n291), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n832), .A2(new_n283), .B1(new_n761), .B2(new_n1007), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n763), .A2(new_n202), .B1(new_n757), .B2(new_n220), .ZN(new_n1033));
  OR4_X1    g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n269), .B1(new_n770), .B2(G326), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n777), .A2(new_n783), .B1(new_n774), .B2(new_n790), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n762), .A2(G317), .B1(G303), .B2(new_n758), .ZN(new_n1037));
  INV_X1    g0837(.A(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n823), .B2(new_n832), .C1(new_n1038), .C2(new_n761), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1035), .B1(new_n526), .B2(new_n766), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1027), .B1(new_n751), .B2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n988), .A2(new_n1016), .B1(new_n1017), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n988), .A2(new_n736), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n686), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n988), .A2(new_n736), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  INV_X1    g0852(.A(new_n686), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1049), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n983), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT110), .ZN(new_n1056));
  MUX2_X1   g0856(.A(new_n981), .B(new_n983), .S(new_n1056), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1057), .B2(new_n1054), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n762), .A2(G311), .B1(new_n760), .B2(G317), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n767), .B2(G107), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n777), .A2(new_n790), .B1(new_n1038), .B2(new_n769), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT114), .Z(new_n1064));
  NOR2_X1   g0864(.A1(new_n774), .A2(new_n526), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n271), .B1(new_n783), .B2(new_n757), .C1(new_n832), .C2(new_n791), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT115), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n763), .A2(new_n1007), .B1(new_n761), .B2(new_n313), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n755), .A2(G50), .B1(new_n347), .B2(new_n758), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1070), .A2(new_n1071), .B1(new_n1073), .B2(KEYINPUT112), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n774), .A2(new_n323), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n271), .B1(new_n770), .B2(G143), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n827), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT112), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1072), .A2(new_n1080), .B1(new_n778), .B2(G68), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1074), .A2(new_n1075), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT115), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n1067), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n751), .B1(new_n1069), .B2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n798), .A2(new_n243), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n802), .B1(new_n492), .B2(new_n210), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n742), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n748), .B2(new_n925), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1057), .B2(new_n1016), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1058), .A2(new_n1090), .ZN(G390));
  NOR2_X1   g0891(.A1(new_n885), .A2(new_n874), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT39), .B1(new_n862), .B2(new_n869), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n874), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n870), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n883), .B1(new_n708), .B2(new_n814), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n881), .B(KEYINPUT116), .Z(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n733), .A2(new_n814), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n881), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1096), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n673), .B1(new_n893), .B2(new_n732), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n895), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1092), .B1(new_n863), .B2(new_n872), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n467), .A2(new_n1106), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n888), .A2(new_n658), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1106), .A2(new_n814), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1100), .A2(new_n1114), .B1(new_n1103), .B2(new_n881), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1103), .B2(new_n881), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n815), .A2(new_n884), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1115), .A2(new_n1099), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1105), .A2(new_n1111), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT117), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT117), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1105), .A2(new_n1111), .A3(new_n1119), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n686), .C1(new_n1125), .C2(new_n1119), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n746), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n742), .B1(new_n820), .B2(new_n347), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT118), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n832), .A2(new_n268), .B1(new_n769), .B2(new_n783), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n763), .A2(new_n526), .B1(new_n757), .B2(new_n492), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n269), .B(new_n1076), .C1(G283), .C2(new_n760), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n778), .A2(G87), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n835), .ZN(new_n1135));
  INV_X1    g0935(.A(G128), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n269), .B1(new_n1007), .B2(new_n774), .C1(new_n761), .C2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n832), .A2(new_n831), .B1(new_n757), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G132), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n763), .A2(new_n1140), .B1(new_n769), .B2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n202), .B2(new_n766), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n778), .A2(G150), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1135), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1129), .B1(new_n1147), .B2(new_n751), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT119), .Z(new_n1149));
  AOI22_X1  g0949(.A1(new_n1125), .A2(new_n1016), .B1(new_n1127), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1126), .A2(new_n1150), .ZN(G378));
  OAI21_X1  g0951(.A(G330), .B1(new_n898), .B2(new_n903), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n343), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n332), .A2(new_n664), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1152), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(G330), .C1(new_n898), .C2(new_n903), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1164), .A2(new_n887), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n887), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1113), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1124), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT122), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1053), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT122), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1113), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n1168), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1163), .A2(new_n746), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n742), .B1(new_n820), .B2(G50), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G33), .A2(G41), .ZN(new_n1181));
  INV_X1    g0981(.A(G41), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G50), .B(new_n1181), .C1(new_n271), .C2(new_n1182), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n763), .A2(new_n1136), .B1(new_n757), .B2(new_n831), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n832), .A2(new_n1140), .B1(new_n761), .B2(new_n1141), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G150), .C2(new_n837), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n777), .B2(new_n1138), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT121), .B(G124), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1181), .B1(new_n769), .B2(new_n1189), .C1(new_n766), .C2(new_n1007), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1187), .B2(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1183), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G41), .B(new_n269), .C1(new_n770), .C2(G283), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n351), .B2(new_n766), .C1(new_n323), .C2(new_n777), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT120), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n763), .A2(new_n268), .B1(new_n291), .B2(new_n757), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n832), .A2(new_n492), .B1(new_n761), .B2(new_n526), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G68), .C2(new_n837), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(KEYINPUT58), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1192), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT58), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1180), .B1(new_n1202), .B2(new_n751), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1178), .A2(new_n1016), .B1(new_n1179), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1177), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1207), .A2(new_n1119), .A3(new_n990), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1100), .A2(new_n746), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n763), .A2(new_n790), .B1(new_n757), .B2(new_n268), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n761), .A2(new_n783), .B1(new_n769), .B2(new_n791), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n271), .B1(new_n832), .B2(new_n526), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1031), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G77), .A2(new_n767), .B1(new_n778), .B2(G97), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n269), .B1(new_n202), .B2(new_n774), .C1(new_n761), .C2(new_n1140), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n763), .A2(new_n831), .B1(new_n757), .B2(new_n313), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n832), .A2(new_n1138), .B1(new_n769), .B2(new_n1136), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G58), .A2(new_n767), .B1(new_n778), .B2(G159), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1213), .A2(new_n1214), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n742), .B1(G68), .B2(new_n820), .C1(new_n1220), .C2(new_n752), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1118), .A2(new_n972), .B1(new_n1209), .B2(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1208), .A2(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G378), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1177), .A2(new_n1224), .A3(new_n1204), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G390), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n1014), .A3(new_n992), .A4(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .ZN(G407));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1119), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1053), .B1(new_n1236), .B2(new_n1207), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1206), .B1(new_n1119), .B2(new_n1235), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1222), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G384), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n844), .B(new_n1222), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G343), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G213), .A3(G2897), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1242), .B(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT125), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1224), .B1(new_n1177), .B2(new_n1204), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1243), .A2(G213), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1204), .A2(new_n1126), .A3(new_n1150), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1175), .A2(new_n990), .A3(new_n1168), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1246), .B(new_n1249), .C1(new_n1250), .C2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(G375), .B2(G378), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1248), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1250), .A2(KEYINPUT62), .A3(new_n1254), .A4(new_n1247), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1227), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n992), .A2(new_n1014), .A3(G390), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(G396), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n992), .A2(new_n1014), .A3(G390), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G390), .B1(new_n992), .B2(new_n1014), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT126), .B(new_n1267), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(KEYINPUT127), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1267), .B1(new_n1265), .B2(KEYINPUT126), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1272), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1250), .A2(new_n1254), .A3(new_n1247), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(KEYINPUT63), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1254), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(new_n1248), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(KEYINPUT124), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1282), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1248), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n1256), .A3(new_n1255), .A4(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1262), .A2(new_n1278), .B1(new_n1287), .B2(new_n1290), .ZN(G405));
  OAI21_X1  g1091(.A(new_n1248), .B1(new_n1226), .B2(new_n1250), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1282), .A2(new_n1225), .A3(new_n1247), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1273), .A2(new_n1277), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


