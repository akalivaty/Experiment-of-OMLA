//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT10), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .A3(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G128), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n204), .A2(KEYINPUT80), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT80), .B1(new_n204), .B2(new_n206), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n207), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT3), .A3(G107), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(G104), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(KEYINPUT3), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n222), .B(KEYINPUT3), .C1(new_n216), .C2(G107), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n220), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n223), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n228), .B2(new_n219), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n197), .B1(new_n215), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n220), .B1(new_n224), .B2(new_n226), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n201), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n203), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT0), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(new_n246), .A3(G101), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n234), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n231), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT65), .B1(new_n251), .B2(G134), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G137), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT11), .B1(new_n254), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n251), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n250), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n250), .A3(new_n260), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT83), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n227), .A2(new_n266), .A3(new_n229), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n227), .B2(new_n229), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n236), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n210), .A2(new_n212), .B1(G143), .B2(new_n201), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n238), .B1(new_n271), .B2(KEYINPUT67), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n274));
  INV_X1    g088(.A(new_n235), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n270), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT10), .B1(new_n277), .B2(new_n214), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n269), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n230), .A2(KEYINPUT81), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n227), .A2(new_n266), .A3(new_n229), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT67), .B(new_n235), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(G128), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n236), .ZN(new_n288));
  INV_X1    g102(.A(new_n214), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n197), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT82), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n249), .B(new_n265), .C1(new_n280), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n288), .A2(new_n289), .A3(new_n230), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n208), .A2(new_n214), .ZN(new_n295));
  INV_X1    g109(.A(new_n207), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n230), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n264), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n299), .A2(KEYINPUT84), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(KEYINPUT84), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n214), .B1(new_n287), .B2(new_n236), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n230), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n230), .B2(new_n215), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(KEYINPUT84), .A3(new_n299), .A4(new_n264), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n196), .B1(new_n293), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n231), .A2(new_n248), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n279), .B1(new_n269), .B2(new_n278), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n283), .A2(KEYINPUT82), .A3(new_n290), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n196), .B1(new_n312), .B2(new_n265), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n249), .B1(new_n280), .B2(new_n291), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n264), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n308), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n192), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n292), .A2(new_n306), .A3(new_n302), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n196), .A2(new_n320), .B1(new_n313), .B2(new_n315), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT85), .B(G469), .C1(new_n321), .C2(G902), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n293), .A2(new_n307), .A3(new_n196), .ZN(new_n324));
  INV_X1    g138(.A(new_n196), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n315), .B2(new_n292), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n318), .B(new_n190), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n264), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n292), .B1(new_n312), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n196), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n302), .A2(new_n306), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n313), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT86), .A3(new_n318), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n191), .B1(new_n323), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G234), .ZN(new_n339));
  OAI21_X1  g153(.A(G217), .B1(new_n339), .B2(G902), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT74), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n187), .A2(new_n339), .A3(G953), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G125), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(G125), .ZN(new_n350));
  INV_X1    g164(.A(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G140), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT16), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT76), .A4(G125), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n201), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n349), .A2(new_n353), .A3(G146), .A4(new_n354), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT24), .B(G110), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n238), .A2(G119), .ZN(new_n361));
  INV_X1    g175(.A(G119), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G128), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n363), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT75), .B1(new_n367), .B2(new_n359), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n362), .A2(G128), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n369), .B(new_n363), .C1(new_n370), .C2(KEYINPUT23), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n366), .A2(new_n368), .B1(G110), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n351), .A2(KEYINPUT16), .A3(G140), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n374), .A2(KEYINPUT16), .B1(new_n375), .B2(KEYINPUT76), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n376), .A2(KEYINPUT77), .A3(G146), .A4(new_n349), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n357), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n201), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n371), .A2(G110), .B1(new_n360), .B2(new_n364), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n373), .A2(new_n382), .A3(KEYINPUT78), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n373), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n344), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(new_n344), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n341), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n388), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n373), .A2(new_n382), .A3(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n396), .B2(new_n344), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT25), .B1(new_n397), .B2(G902), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n341), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G902), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n392), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n362), .A2(G116), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT69), .B(G116), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(G119), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT2), .B(G113), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(KEYINPUT68), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(KEYINPUT68), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n251), .A2(G134), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n254), .A2(G137), .ZN(new_n417));
  OAI21_X1  g231(.A(G131), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n263), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n288), .B2(new_n289), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n244), .B1(new_n262), .B2(new_n263), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n414), .B(new_n415), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n263), .A2(new_n418), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n277), .B2(new_n214), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n256), .A2(new_n250), .A3(new_n260), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n245), .B1(new_n425), .B2(new_n261), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n424), .A2(KEYINPUT68), .A3(new_n413), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n412), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G237), .A2(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G210), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT27), .Z(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT26), .B(G101), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n426), .B(new_n412), .C1(new_n303), .C2(new_n419), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR4_X1   g249(.A1(new_n428), .A2(KEYINPUT31), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT71), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n412), .B1(new_n424), .B2(new_n426), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT72), .B1(new_n435), .B2(KEYINPUT28), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n436), .A2(new_n437), .B1(new_n433), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n422), .A2(new_n427), .ZN(new_n446));
  INV_X1    g260(.A(new_n411), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n410), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT31), .ZN(new_n450));
  INV_X1    g264(.A(new_n433), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .A4(new_n434), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT71), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n428), .A2(new_n433), .A3(new_n435), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n451), .A3(new_n434), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n445), .A2(new_n453), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(G472), .A2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND4_X1   g277(.A1(new_n451), .A2(new_n439), .A3(new_n440), .A4(new_n443), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n464), .B2(KEYINPUT29), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n433), .B1(new_n428), .B2(new_n435), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n439), .A2(new_n440), .A3(new_n451), .A4(new_n443), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n459), .A2(new_n463), .B1(new_n472), .B2(G472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n455), .A2(new_n437), .A3(new_n450), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n444), .A2(new_n433), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n453), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n456), .A2(new_n458), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n460), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n407), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n234), .A2(new_n448), .A3(new_n247), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n234), .A2(KEYINPUT87), .A3(new_n448), .A4(new_n247), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n488));
  INV_X1    g302(.A(G113), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT5), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n408), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n488), .A2(new_n491), .B1(new_n410), .B2(new_n447), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n267), .B2(new_n268), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n483), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n484), .A2(new_n485), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(new_n482), .A3(new_n493), .A4(new_n487), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n303), .A2(new_n351), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n244), .A2(G125), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n194), .A2(G224), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n501), .B(new_n502), .Z(new_n503));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n504), .B(new_n483), .C1(new_n486), .C2(new_n494), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(G224), .A3(new_n194), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n499), .A2(KEYINPUT7), .A3(new_n502), .A4(new_n500), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n492), .A2(new_n230), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n492), .A2(new_n230), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n482), .B(KEYINPUT8), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AND4_X1   g328(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n515), .B2(new_n497), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n506), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n517), .B(KEYINPUT88), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n506), .B2(new_n516), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n481), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n506), .A2(new_n516), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n520), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n518), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n481), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n350), .A2(new_n352), .A3(new_n201), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n201), .B1(new_n350), .B2(new_n352), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT91), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n350), .A2(new_n352), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G146), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n380), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT18), .A2(G131), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n199), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(G214), .B2(new_n429), .ZN(new_n542));
  INV_X1    g356(.A(G237), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n194), .A3(G214), .ZN(new_n544));
  NOR2_X1   g358(.A1(KEYINPUT90), .A2(G143), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n539), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(G214), .A3(new_n429), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT18), .A4(G131), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n534), .A2(new_n538), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n357), .B(KEYINPUT77), .ZN(new_n552));
  OAI21_X1  g366(.A(G131), .B1(new_n542), .B2(new_n546), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n549), .A3(new_n250), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n535), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n374), .A2(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n553), .A2(new_n554), .B1(new_n558), .B2(new_n201), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n551), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G113), .B(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(new_n216), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT92), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n538), .A2(new_n534), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n547), .A2(new_n550), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n553), .A2(new_n554), .ZN(new_n567));
  INV_X1    g381(.A(new_n558), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(G146), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n377), .A2(new_n379), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n572));
  INV_X1    g386(.A(new_n562), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(new_n567), .B2(KEYINPUT17), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n553), .A2(new_n576), .A3(new_n577), .A4(new_n554), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT17), .B(G131), .C1(new_n542), .C2(new_n546), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n356), .A2(new_n357), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n562), .A3(new_n566), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n563), .A2(new_n574), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G475), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n531), .B1(new_n585), .B2(KEYINPUT20), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT20), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT94), .B(new_n587), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n587), .A3(new_n584), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n409), .A2(KEYINPUT14), .A3(G122), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n409), .A2(G122), .ZN(new_n593));
  INV_X1    g407(.A(G122), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G116), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(G107), .B(new_n592), .C1(new_n596), .C2(KEYINPUT14), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n199), .A2(G128), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n238), .A2(G143), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G134), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n599), .A3(new_n254), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(KEYINPUT97), .A3(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n593), .B2(new_n595), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n593), .A2(new_n608), .A3(new_n595), .ZN(new_n611));
  AOI21_X1  g425(.A(G107), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n599), .B1(new_n598), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n598), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT96), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n598), .A2(new_n619), .A3(new_n615), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n602), .B1(new_n621), .B2(new_n254), .ZN(new_n622));
  INV_X1    g436(.A(new_n611), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n218), .B1(new_n623), .B2(new_n609), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n610), .A2(G107), .A3(new_n611), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G217), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n188), .A2(new_n628), .A3(G953), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n614), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n629), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n613), .B2(new_n626), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G478), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(KEYINPUT15), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n581), .A2(new_n566), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n573), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n582), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n190), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(G475), .ZN(new_n642));
  INV_X1    g456(.A(G952), .ZN(new_n643));
  AOI211_X1 g457(.A(G953), .B(new_n643), .C1(G234), .C2(G237), .ZN(new_n644));
  OAI211_X1 g458(.A(G902), .B(G953), .C1(new_n339), .C2(new_n543), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT21), .B(G898), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n591), .A2(new_n637), .A3(new_n642), .A4(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n338), .A2(new_n480), .A3(new_n530), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT99), .B(G101), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G3));
  INV_X1    g466(.A(G472), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n459), .B2(new_n190), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n453), .A2(new_n474), .A3(new_n475), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n456), .A2(new_n458), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n461), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n338), .A2(new_n406), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n648), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n517), .B1(new_n506), .B2(new_n516), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n481), .B(new_n660), .C1(new_n519), .C2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n630), .A2(new_n632), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT33), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT33), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n630), .A2(new_n632), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(G478), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n634), .A2(new_n190), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n633), .B2(new_n634), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT94), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n585), .A2(new_n531), .A3(KEYINPUT20), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n589), .ZN(new_n675));
  INV_X1    g489(.A(new_n642), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n663), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n659), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT34), .B(G104), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  INV_X1    g495(.A(new_n191), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT86), .B1(new_n335), .B2(new_n318), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n331), .A2(new_n196), .B1(new_n313), .B2(new_n333), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n684), .A2(new_n328), .A3(G469), .A4(G902), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n319), .A2(new_n322), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n476), .A2(new_n477), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n478), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n688), .A2(new_n407), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n636), .A2(new_n642), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n673), .A2(new_n694), .A3(new_n674), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT100), .B1(new_n586), .B2(new_n588), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT101), .B1(new_n697), .B2(new_n589), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n699), .B(new_n590), .C1(new_n695), .C2(new_n696), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n663), .B(new_n693), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(KEYINPUT102), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(KEYINPUT102), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n692), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT35), .B(G107), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G9));
  OAI211_X1 g520(.A(new_n394), .B(new_n395), .C1(KEYINPUT36), .C2(new_n344), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n344), .A2(KEYINPUT36), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n383), .B2(new_n384), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n707), .A2(new_n402), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n400), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n654), .A2(new_n657), .A3(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n338), .A2(new_n530), .A3(new_n649), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT37), .B(G110), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G12));
  INV_X1    g529(.A(G900), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n646), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  INV_X1    g532(.A(new_n644), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n693), .B(new_n722), .C1(new_n698), .C2(new_n700), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n481), .B1(new_n519), .B2(new_n661), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n711), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n472), .A2(G472), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT32), .B1(new_n459), .B2(new_n460), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n688), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G128), .ZN(G30));
  OAI21_X1  g548(.A(new_n451), .B1(new_n428), .B2(new_n435), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n435), .A2(new_n438), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n735), .B(new_n190), .C1(new_n451), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G472), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n479), .A2(new_n728), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT104), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n722), .B(KEYINPUT39), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n338), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(KEYINPUT40), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(KEYINPUT40), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n527), .B(KEYINPUT38), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n636), .B1(new_n675), .B2(new_n676), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n481), .A3(new_n711), .A4(new_n746), .ZN(new_n747));
  OR4_X1    g561(.A1(new_n740), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  INV_X1    g563(.A(new_n671), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(new_n722), .C1(new_n591), .C2(new_n642), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT105), .B1(new_n751), .B2(new_n724), .ZN(new_n752));
  INV_X1    g566(.A(new_n481), .ZN(new_n753));
  INV_X1    g567(.A(new_n517), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n525), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n755), .B2(new_n518), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n677), .A3(new_n757), .A4(new_n722), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n711), .B1(new_n473), .B2(new_n479), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n338), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G146), .ZN(G48));
  OAI21_X1  g576(.A(new_n406), .B1(new_n729), .B2(new_n730), .ZN(new_n763));
  OAI21_X1  g577(.A(G469), .B1(new_n684), .B2(G902), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n337), .A2(new_n682), .A3(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n678), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT41), .B(G113), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G15));
  INV_X1    g582(.A(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n480), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n702), .B2(new_n703), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  NAND4_X1  g587(.A1(new_n337), .A2(new_n682), .A3(new_n756), .A4(new_n764), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n649), .A3(new_n760), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G119), .ZN(G21));
  AOI21_X1  g591(.A(KEYINPUT106), .B1(new_n399), .B2(new_n404), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n779), .B(new_n405), .C1(new_n391), .C2(new_n398), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n457), .A2(KEYINPUT31), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n461), .B1(new_n655), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n654), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n637), .B1(new_n591), .B2(new_n642), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n724), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n769), .A2(new_n784), .A3(new_n660), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G122), .ZN(G24));
  INV_X1    g602(.A(new_n722), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n671), .C1(new_n675), .C2(new_n676), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n655), .A2(new_n782), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n460), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n690), .A2(new_n790), .A3(new_n726), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n774), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n351), .ZN(G27));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n526), .A2(new_n481), .A3(new_n518), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n191), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT107), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n308), .A2(new_n316), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n318), .B1(new_n800), .B2(new_n190), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n337), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(KEYINPUT107), .B(new_n801), .C1(new_n329), .C2(new_n336), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n480), .B(new_n798), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n796), .B1(new_n805), .B2(new_n751), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n729), .B1(KEYINPUT108), .B2(new_n479), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n479), .A2(KEYINPUT108), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n781), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n798), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n802), .B1(new_n683), .B2(new_n685), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT107), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n337), .A2(new_n799), .A3(new_n802), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n751), .A2(new_n796), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G131), .ZN(G33));
  INV_X1    g632(.A(new_n723), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n819), .A3(new_n480), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  NAND2_X1  g635(.A1(new_n691), .A2(new_n726), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT109), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n586), .A2(new_n588), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n642), .B1(new_n824), .B2(new_n589), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n750), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT43), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT44), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n797), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n823), .A2(KEYINPUT44), .A3(new_n828), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT45), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n800), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n321), .A2(KEYINPUT45), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(G469), .ZN(new_n837));
  NAND2_X1  g651(.A1(G469), .A2(G902), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT46), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n337), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n682), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n741), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(KEYINPUT110), .B(G137), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(G39));
  INV_X1    g663(.A(KEYINPUT47), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n790), .A2(new_n832), .A3(new_n407), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n730), .A3(new_n729), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT111), .B(G140), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(G42));
  NAND2_X1  g672(.A1(new_n337), .A2(new_n764), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT49), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n682), .A2(new_n481), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n745), .A2(new_n781), .A3(new_n826), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n740), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n650), .A2(new_n713), .A3(new_n776), .A4(new_n787), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT112), .B1(new_n825), .B2(new_n671), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n677), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n825), .B2(new_n637), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n591), .A2(KEYINPUT113), .A3(new_n636), .A4(new_n642), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n866), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n648), .B1(new_n524), .B2(new_n529), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n659), .A2(new_n874), .B1(new_n770), .B2(new_n678), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n697), .A2(new_n589), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n699), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n697), .A2(KEYINPUT101), .A3(new_n589), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n797), .A2(new_n642), .A3(new_n637), .A4(new_n789), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n732), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n793), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n814), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n820), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n876), .A2(new_n885), .A3(new_n772), .A4(new_n817), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n654), .A2(new_n783), .A3(new_n711), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n775), .A2(new_n790), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n880), .A2(new_n756), .A3(new_n693), .A4(new_n722), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n338), .A2(new_n760), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n710), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n722), .B(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n190), .B1(new_n403), .B2(new_n392), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n401), .B1(new_n896), .B2(KEYINPUT25), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n389), .A2(new_n390), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n892), .B(new_n895), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n399), .A2(KEYINPUT115), .A3(new_n892), .A4(new_n895), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n682), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n785), .A3(new_n724), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n739), .B(new_n904), .C1(new_n803), .C2(new_n804), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n761), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT52), .B1(new_n891), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n794), .B1(new_n725), .B2(new_n732), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n812), .A2(new_n813), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n728), .A2(new_n738), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n730), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n710), .B(new_n894), .C1(new_n391), .C2(new_n398), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n191), .B1(new_n912), .B2(KEYINPUT115), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n756), .A3(new_n746), .A4(new_n901), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n732), .A2(new_n759), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT52), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n864), .B1(new_n886), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n907), .A2(new_n918), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n872), .A2(new_n873), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n766), .B1(new_n922), .B2(new_n692), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n650), .A2(new_n713), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n776), .A2(new_n787), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n772), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n820), .A2(new_n882), .A3(new_n884), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n806), .B2(new_n816), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n921), .A2(new_n926), .A3(new_n928), .A4(KEYINPUT53), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n920), .A2(new_n929), .A3(KEYINPUT54), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n828), .A2(new_n644), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n769), .A2(new_n832), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(KEYINPUT118), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n809), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n943), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n936), .A2(new_n407), .A3(new_n719), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n677), .A3(new_n740), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n828), .A2(new_n644), .A3(new_n784), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n643), .B(G953), .C1(new_n947), .C2(new_n775), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n946), .B(new_n948), .C1(new_n943), .C2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT51), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n745), .A2(new_n765), .A3(new_n481), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT117), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n945), .A2(new_n825), .A3(new_n671), .A4(new_n740), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n887), .B1(new_n938), .B2(new_n940), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n947), .A2(new_n832), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n859), .A2(new_n682), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n853), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n957), .A2(new_n958), .A3(new_n952), .A4(new_n959), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT116), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n853), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n851), .A2(KEYINPUT116), .A3(new_n852), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n967), .B(new_n968), .C1(new_n682), .C2(new_n859), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n965), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n951), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n934), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(G952), .A2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n863), .B1(new_n972), .B2(new_n973), .ZN(G75));
  NOR2_X1   g788(.A1(new_n194), .A2(G952), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n190), .B1(new_n920), .B2(new_n929), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT56), .B1(new_n977), .B2(G210), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n498), .A2(new_n505), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n503), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT121), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n976), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT122), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n930), .B2(G902), .ZN(new_n986));
  AOI211_X1 g800(.A(KEYINPUT122), .B(new_n190), .C1(new_n920), .C2(new_n929), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n520), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT56), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n989), .B2(new_n991), .ZN(G51));
  INV_X1    g806(.A(new_n837), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n838), .B(KEYINPUT57), .Z(new_n995));
  NAND3_X1  g809(.A1(new_n932), .A2(new_n933), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n326), .B2(new_n324), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n975), .B1(new_n994), .B2(new_n997), .ZN(G54));
  AND2_X1   g812(.A1(KEYINPUT58), .A2(G475), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n583), .B1(new_n988), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n805), .ZN(new_n1001));
  AOI22_X1  g815(.A1(new_n1001), .A2(new_n819), .B1(new_n883), .B2(new_n814), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n817), .A2(new_n1002), .A3(new_n882), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n772), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT53), .B1(new_n1005), .B2(new_n921), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n886), .A2(new_n864), .A3(new_n919), .ZN(new_n1007));
  OAI21_X1  g821(.A(G902), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(KEYINPUT122), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n977), .A2(new_n985), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n583), .A2(new_n999), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n976), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1000), .A2(new_n1013), .ZN(G60));
  NAND2_X1  g828(.A1(new_n665), .A2(new_n667), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n669), .B(KEYINPUT59), .Z(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n934), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n932), .A2(new_n1015), .A3(new_n933), .A4(new_n1016), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n976), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1017), .A2(new_n1019), .ZN(G63));
  XNOR2_X1  g834(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n628), .A2(new_n190), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n930), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n397), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n930), .A2(new_n709), .A3(new_n707), .A4(new_n1023), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1025), .A2(new_n976), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT61), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1025), .A2(KEYINPUT61), .A3(new_n976), .A4(new_n1026), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(G66));
  INV_X1    g845(.A(G224), .ZN(new_n1032));
  OAI21_X1  g846(.A(G953), .B1(new_n647), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n926), .B2(G953), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n979), .B1(G898), .B2(new_n194), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT124), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1034), .B(new_n1036), .ZN(G69));
  XNOR2_X1  g851(.A(new_n446), .B(new_n568), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n742), .A2(new_n797), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1039), .A2(new_n480), .A3(new_n872), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n847), .A2(new_n856), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n908), .A2(new_n761), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n908), .A2(KEYINPUT125), .A3(new_n761), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n748), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT62), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g862(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1049), .A2(KEYINPUT62), .A3(new_n748), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1041), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1038), .B1(new_n1051), .B2(G953), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1038), .B1(G900), .B2(G953), .ZN(new_n1053));
  AOI22_X1  g867(.A1(new_n853), .A2(new_n855), .B1(new_n819), .B2(new_n1001), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n846), .A2(new_n786), .A3(new_n809), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n1056), .A2(new_n817), .A3(new_n847), .A4(new_n1049), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1053), .B1(new_n1057), .B2(G953), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1060), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1052), .A2(new_n1062), .A3(new_n1058), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1061), .A2(new_n1063), .ZN(G72));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  NAND2_X1  g880(.A1(new_n457), .A2(new_n467), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n930), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g882(.A(new_n1066), .B(KEYINPUT126), .Z(new_n1069));
  AOI21_X1  g883(.A(new_n1069), .B1(new_n1051), .B2(new_n926), .ZN(new_n1070));
  OAI211_X1 g884(.A(new_n976), .B(new_n1068), .C1(new_n1070), .C2(new_n735), .ZN(new_n1071));
  NAND3_X1  g885(.A1(new_n449), .A2(new_n433), .A3(new_n434), .ZN(new_n1072));
  NAND4_X1  g886(.A1(new_n847), .A2(new_n1054), .A3(new_n817), .A4(new_n1055), .ZN(new_n1073));
  INV_X1    g887(.A(new_n1049), .ZN(new_n1074));
  NOR3_X1   g888(.A1(new_n1073), .A2(new_n1004), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g889(.A(KEYINPUT127), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT127), .ZN(new_n1077));
  INV_X1    g891(.A(new_n1069), .ZN(new_n1078));
  OAI211_X1 g892(.A(new_n1077), .B(new_n1078), .C1(new_n1057), .C2(new_n1004), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1072), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g894(.A1(new_n1071), .A2(new_n1080), .ZN(G57));
endmodule


