//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n444, new_n449, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT69), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT70), .Z(G217));
  NOR4_X1   g029(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g032(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT71), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n459), .A2(G567), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(KEYINPUT72), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n457), .B2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(KEYINPUT72), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT73), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n469), .A2(new_n471), .A3(new_n478), .A4(G125), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n474), .B1(new_n480), .B2(G2105), .ZN(G160));
  NAND2_X1  g056(.A1(new_n469), .A2(new_n471), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n482), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n469), .A2(new_n471), .A3(G126), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT74), .A2(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(G2104), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n483), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n469), .A2(new_n471), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n483), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n498), .A2(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT4), .A4(G138), .ZN(new_n504));
  NAND2_X1  g079(.A1(G102), .A2(G2104), .ZN(new_n505));
  AOI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AND3_X1   g090(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(new_n510), .B2(new_n511), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n519), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n530), .B(new_n531), .C1(new_n513), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n518), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT76), .B(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n513), .A2(new_n537), .B1(new_n518), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(G171));
  XOR2_X1   g117(.A(KEYINPUT77), .B(G43), .Z(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n513), .A2(new_n543), .B1(new_n544), .B2(new_n518), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n526), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NOR2_X1   g129(.A1(new_n516), .A2(new_n517), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(new_n558), .A3(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n526), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n534), .A2(G91), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n510), .A2(new_n511), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n521), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  OR2_X1    g149(.A1(new_n519), .A2(new_n527), .ZN(G303));
  NAND3_X1  g150(.A1(new_n512), .A2(G49), .A3(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n565), .A2(new_n578), .A3(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n534), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(G288));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n518), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n555), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n524), .A2(KEYINPUT81), .A3(G61), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n585), .B1(new_n591), .B2(G651), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n513), .A2(new_n594), .B1(new_n595), .B2(new_n518), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n526), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n557), .A2(new_n558), .A3(G66), .ZN(new_n602));
  INV_X1    g177(.A(G79), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n521), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(G651), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n565), .A2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n534), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  NAND3_X1  g186(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n484), .A2(G123), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT83), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n486), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n483), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT84), .B(G2096), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT12), .B1(new_n501), .B2(new_n468), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n486), .A2(new_n635), .A3(G2104), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  INV_X1    g218(.A(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(KEYINPUT86), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n645), .A2(new_n646), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n650), .A2(KEYINPUT86), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n647), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n642), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(new_n642), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(new_n656), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n641), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  AOI211_X1 g247(.A(KEYINPUT88), .B(new_n672), .C1(new_n666), .C2(new_n667), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n672), .A3(new_n667), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G14), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2067), .B(G2678), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT17), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(new_n692), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n692), .A3(new_n695), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT91), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(G166), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G22), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G23), .ZN(new_n716));
  INV_X1    g291(.A(G288), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT33), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(new_n714), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n711), .A2(G6), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n592), .B2(new_n711), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n715), .A2(new_n720), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT34), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n711), .A2(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n599), .B2(new_n711), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G1986), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(G1986), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n484), .A2(G119), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n486), .A2(G131), .ZN(new_n735));
  OR2_X1    g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n736), .B(G2104), .C1(G107), .C2(new_n483), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n732), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT35), .B(G1991), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT92), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n727), .A2(new_n730), .A3(new_n731), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT36), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n711), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n548), .B2(new_n711), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1341), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n732), .A2(G26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n486), .A2(G140), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n483), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(new_n732), .ZN(new_n756));
  MUX2_X1   g331(.A(new_n749), .B(new_n756), .S(KEYINPUT28), .Z(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n711), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n613), .B2(new_n711), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n748), .B(new_n759), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n486), .A2(G139), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n500), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n770), .C1(new_n483), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G29), .B2(G33), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n711), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n711), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT31), .B(G11), .Z(new_n782));
  OR3_X1    g357(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n732), .A2(G35), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G162), .B2(new_n732), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT29), .B(G2090), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n775), .A2(new_n776), .ZN(new_n788));
  AND2_X1   g363(.A1(KEYINPUT30), .A2(G28), .ZN(new_n789));
  NOR2_X1   g364(.A1(KEYINPUT30), .A2(G28), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n732), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G5), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G171), .B2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n793), .B2(G1961), .ZN(new_n794));
  INV_X1    g369(.A(new_n793), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n794), .B1(new_n797), .B2(KEYINPUT99), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(KEYINPUT99), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n780), .A2(G1966), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n788), .A2(new_n798), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n732), .A2(G27), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G164), .B2(new_n732), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2078), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n783), .A2(new_n787), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n711), .A2(KEYINPUT23), .A3(G20), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n808));
  INV_X1    g383(.A(G20), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n810), .C1(new_n617), .C2(new_n711), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n766), .A2(new_n805), .A3(new_n806), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G29), .A2(G32), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n500), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G129), .B2(new_n484), .ZN(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT26), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n815), .B1(new_n823), .B2(G29), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT27), .B(G1996), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n827));
  NOR2_X1   g402(.A1(KEYINPUT24), .A2(G34), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(KEYINPUT24), .A2(G34), .ZN(new_n830));
  AOI21_X1  g405(.A(G29), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(G160), .A2(G29), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n827), .B2(new_n831), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT97), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G2084), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n745), .A2(new_n814), .A3(new_n826), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n631), .A2(new_n732), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  AOI22_X1  g414(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT100), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G651), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n534), .A2(G93), .B1(new_n565), .B2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT101), .B(G860), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  INV_X1    g422(.A(new_n548), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n844), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n620), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n847), .B1(new_n853), .B2(new_n845), .ZN(G145));
  XNOR2_X1  g429(.A(new_n508), .B(new_n754), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n773), .A2(new_n822), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n773), .A2(new_n822), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n855), .A3(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n500), .A2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n486), .A2(G142), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n483), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n484), .A2(KEYINPUT102), .A3(G130), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n867), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n637), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n739), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n739), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n863), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  INV_X1    g453(.A(new_n874), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(KEYINPUT103), .A3(new_n874), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n860), .A2(new_n862), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n631), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n863), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n882), .ZN(new_n890));
  INV_X1    g465(.A(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n877), .A2(new_n893), .A3(new_n882), .A4(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n887), .A2(new_n892), .A3(new_n897), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(G299), .A2(KEYINPUT106), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n570), .A2(new_n902), .A3(new_n571), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n903), .A3(new_n613), .ZN(new_n904));
  NAND3_X1  g479(.A1(G299), .A2(new_n612), .A3(KEYINPUT106), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n622), .B(new_n849), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(new_n599), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n717), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n717), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n592), .B(KEYINPUT107), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(KEYINPUT108), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n904), .A2(new_n905), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n927));
  AND4_X1   g502(.A1(new_n911), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n911), .A2(new_n926), .B1(new_n924), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n844), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(G868), .B2(new_n931), .ZN(G295));
  OAI21_X1  g507(.A(new_n930), .B1(G868), .B2(new_n931), .ZN(G331));
  NOR2_X1   g508(.A1(G168), .A2(KEYINPUT109), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n849), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n931), .A2(new_n848), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n844), .A2(new_n548), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G301), .B1(KEYINPUT109), .B2(G168), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n941), .B(new_n944), .C1(new_n907), .C2(new_n908), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n925), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n923), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n945), .A2(new_n922), .A3(new_n947), .A4(new_n921), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n949), .A2(new_n951), .A3(new_n954), .A4(new_n950), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G397));
  XOR2_X1   g535(.A(KEYINPUT58), .B(G1341), .Z(new_n961));
  INV_X1    g536(.A(KEYINPUT120), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n480), .A2(G2105), .ZN(new_n963));
  INV_X1    g538(.A(new_n474), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT110), .B(G40), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(G160), .A2(KEYINPUT111), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n482), .A2(new_n502), .A3(G2105), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n469), .A2(new_n471), .A3(G126), .ZN(new_n975));
  AND2_X1   g550(.A1(KEYINPUT74), .A2(G114), .ZN(new_n976));
  NOR2_X1   g551(.A1(KEYINPUT74), .A2(G114), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n468), .ZN(new_n978));
  OAI21_X1  g553(.A(G2105), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n979), .B2(KEYINPUT4), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n973), .B1(new_n980), .B2(new_n506), .ZN(new_n981));
  AOI211_X1 g556(.A(KEYINPUT120), .B(new_n981), .C1(new_n968), .C2(new_n969), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n961), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n985), .A2(new_n986), .B1(new_n968), .B2(new_n969), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n508), .B2(new_n973), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n984), .B(G1384), .C1(new_n503), .C2(new_n507), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT113), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT59), .B1(new_n993), .B2(new_n548), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT59), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n848), .C1(new_n983), .C2(new_n992), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT60), .ZN(new_n998));
  AND4_X1   g573(.A1(KEYINPUT111), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT111), .B1(G160), .B2(new_n965), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n971), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT120), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n970), .A2(new_n962), .A3(new_n971), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n758), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n971), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n970), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n762), .ZN(new_n1010));
  AND4_X1   g585(.A1(new_n998), .A2(new_n1004), .A3(new_n613), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n985), .A2(new_n986), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT56), .B(G2072), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n991), .A2(new_n970), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n999), .A2(new_n1000), .B1(new_n971), .B2(new_n1006), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n812), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT9), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n566), .B(new_n1019), .ZN(new_n1020));
  NOR4_X1   g595(.A1(new_n1020), .A2(new_n561), .A3(KEYINPUT57), .A4(new_n562), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n563), .B2(new_n567), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1014), .A2(new_n1024), .A3(new_n1017), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT61), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1011), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT121), .B(new_n1024), .C1(new_n1014), .C2(new_n1017), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT61), .B(new_n1027), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n998), .B1(new_n1035), .B2(new_n612), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n612), .B2(new_n1035), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n997), .A2(new_n1030), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n613), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1027), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n577), .A2(new_n579), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n580), .A2(new_n581), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(G1976), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(G288), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1001), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n591), .A2(G651), .ZN(new_n1053));
  INV_X1    g628(.A(new_n585), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT116), .B(G1981), .Z(new_n1056));
  AOI211_X1 g631(.A(new_n585), .B(new_n1056), .C1(new_n591), .C2(G651), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1056), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1053), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(new_n1061), .C1(new_n1052), .C2(new_n592), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(G8), .A3(new_n1001), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1001), .A2(G8), .A3(new_n1049), .A4(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1051), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT55), .Z(new_n1069));
  AOI21_X1  g644(.A(G1971), .B1(new_n987), .B2(new_n991), .ZN(new_n1070));
  INV_X1    g645(.A(G2090), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1071), .A2(new_n970), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1072));
  OAI211_X1 g647(.A(G8), .B(new_n1069), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n986), .B1(new_n985), .B2(new_n1076), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n989), .A2(KEYINPUT113), .B1(new_n999), .B2(new_n1000), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n714), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1016), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n981), .A2(new_n1005), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n970), .A3(new_n1071), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1075), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n1069), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1074), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G2078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n987), .A2(new_n1086), .A3(new_n991), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n1088), .B1(new_n796), .B2(new_n1009), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n985), .A2(new_n1076), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1090), .A2(new_n883), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G171), .B(KEYINPUT54), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n989), .A2(new_n990), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n1086), .A3(new_n970), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1098), .A2(KEYINPUT124), .A3(new_n1086), .A4(new_n970), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT53), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1095), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT119), .B(G2084), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n970), .A2(new_n1007), .A3(new_n1008), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1966), .B1(new_n1098), .B2(new_n970), .ZN(new_n1110));
  OAI21_X1  g685(.A(G8), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G286), .A2(G8), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT122), .Z(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1966), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n999), .A2(new_n1000), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1090), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1075), .B1(new_n1120), .B2(new_n1108), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(KEYINPUT51), .A3(new_n1108), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1113), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1117), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1085), .A2(new_n1097), .A3(new_n1106), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1042), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G288), .A2(G1976), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT118), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1060), .B1(new_n1063), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(G8), .A3(new_n1001), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1051), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT117), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1051), .A2(new_n1064), .A3(new_n1137), .A4(new_n1066), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1139), .B2(new_n1073), .ZN(new_n1140));
  OAI21_X1  g715(.A(G8), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1069), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT63), .A3(new_n1073), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1111), .A2(G286), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1144), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1067), .B(new_n1073), .C1(new_n1069), .C2(new_n1083), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1140), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1129), .A2(new_n1130), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1127), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1140), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n1085), .B2(new_n1145), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1144), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT126), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n1149), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1160), .A2(G171), .A3(new_n1104), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1152), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n970), .A2(new_n989), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n988), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n822), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT112), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n754), .B(new_n758), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n823), .B2(new_n988), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n741), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n738), .B(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n599), .B(G1986), .Z(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1165), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1163), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n739), .A3(new_n1172), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n755), .A2(new_n758), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1164), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OR3_X1    g755(.A1(new_n1164), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  NOR2_X1   g757(.A1(new_n1174), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT46), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT127), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1166), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1169), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1165), .B1(new_n822), .B2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1186), .B(new_n1188), .C1(KEYINPUT127), .C2(new_n1184), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT47), .Z(new_n1190));
  NOR3_X1   g765(.A1(new_n1180), .A2(new_n1183), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g767(.A(new_n466), .B(G401), .C1(new_n896), .C2(new_n898), .ZN(new_n1194));
  NOR2_X1   g768(.A1(G229), .A2(G227), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n1194), .A2(new_n1195), .A3(new_n956), .ZN(G308));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(new_n956), .ZN(G225));
endmodule


