

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739;

  AND2_X1 U374 ( .A1(n528), .A2(n414), .ZN(n529) );
  NOR2_X1 U375 ( .A1(G902), .A2(n693), .ZN(n499) );
  XNOR2_X1 U376 ( .A(n449), .B(n448), .ZN(n496) );
  XOR2_X1 U377 ( .A(KEYINPUT68), .B(KEYINPUT4), .Z(n351) );
  XNOR2_X2 U378 ( .A(n512), .B(n511), .ZN(n376) );
  INV_X1 U379 ( .A(G953), .ZN(n726) );
  XNOR2_X2 U380 ( .A(n439), .B(G472), .ZN(n657) );
  NAND2_X2 U381 ( .A1(n552), .A2(n457), .ZN(n404) );
  XNOR2_X2 U382 ( .A(n452), .B(KEYINPUT19), .ZN(n552) );
  NOR2_X2 U383 ( .A1(n376), .A2(n513), .ZN(n514) );
  NOR2_X1 U384 ( .A1(n653), .A2(n500), .ZN(n650) );
  XNOR2_X1 U385 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n441) );
  NAND2_X1 U386 ( .A1(n529), .A2(n530), .ZN(n532) );
  XNOR2_X1 U387 ( .A(n425), .B(n424), .ZN(n653) );
  NAND2_X1 U388 ( .A1(n429), .A2(n428), .ZN(n478) );
  XNOR2_X1 U389 ( .A(n399), .B(G125), .ZN(n442) );
  XNOR2_X1 U390 ( .A(n381), .B(n380), .ZN(n597) );
  NOR2_X1 U391 ( .A1(n724), .A2(n597), .ZN(n385) );
  XOR2_X1 U392 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n466) );
  XNOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n465) );
  XOR2_X1 U394 ( .A(G122), .B(G104), .Z(n464) );
  NAND2_X1 U395 ( .A1(n586), .A2(n396), .ZN(n395) );
  AND2_X1 U396 ( .A1(n352), .A2(n587), .ZN(n396) );
  NOR2_X1 U397 ( .A1(n738), .A2(n508), .ZN(n509) );
  NOR2_X1 U398 ( .A1(n373), .A2(n370), .ZN(n508) );
  NAND2_X1 U399 ( .A1(n374), .A2(n559), .ZN(n373) );
  XNOR2_X1 U400 ( .A(n442), .B(n398), .ZN(n461) );
  INV_X1 U401 ( .A(KEYINPUT10), .ZN(n398) );
  XNOR2_X1 U402 ( .A(G131), .B(G134), .ZN(n718) );
  AND2_X1 U403 ( .A1(n566), .A2(n541), .ZN(n402) );
  INV_X1 U404 ( .A(n549), .ZN(n403) );
  OR2_X1 U405 ( .A1(G237), .A2(G902), .ZN(n451) );
  INV_X1 U406 ( .A(KEYINPUT30), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n418), .B(n367), .ZN(n479) );
  INV_X1 U408 ( .A(KEYINPUT8), .ZN(n367) );
  XNOR2_X1 U409 ( .A(G128), .B(G119), .ZN(n415) );
  XOR2_X1 U410 ( .A(KEYINPUT24), .B(G110), .Z(n416) );
  XNOR2_X1 U411 ( .A(n461), .B(n397), .ZN(n717) );
  INV_X1 U412 ( .A(n493), .ZN(n397) );
  XOR2_X1 U413 ( .A(G137), .B(G140), .Z(n493) );
  NAND2_X1 U414 ( .A1(n601), .A2(n600), .ZN(n616) );
  XNOR2_X1 U415 ( .A(n545), .B(KEYINPUT39), .ZN(n576) );
  XNOR2_X1 U416 ( .A(n357), .B(n355), .ZN(n520) );
  INV_X1 U417 ( .A(n590), .ZN(n407) );
  NOR2_X2 U418 ( .A1(n520), .A2(n570), .ZN(n523) );
  NAND2_X1 U419 ( .A1(n616), .A2(n412), .ZN(n413) );
  AND2_X1 U420 ( .A1(n615), .A2(G210), .ZN(n412) );
  INV_X1 U421 ( .A(KEYINPUT90), .ZN(n375) );
  INV_X1 U422 ( .A(G146), .ZN(n399) );
  NAND2_X1 U423 ( .A1(G953), .A2(G902), .ZN(n535) );
  XNOR2_X1 U424 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n432) );
  XOR2_X1 U425 ( .A(G137), .B(KEYINPUT88), .Z(n433) );
  XNOR2_X1 U426 ( .A(n410), .B(n431), .ZN(n440) );
  XNOR2_X1 U427 ( .A(G113), .B(G116), .ZN(n431) );
  XNOR2_X1 U428 ( .A(n411), .B(G119), .ZN(n410) );
  INV_X1 U429 ( .A(KEYINPUT3), .ZN(n411) );
  XOR2_X1 U430 ( .A(KEYINPUT9), .B(G122), .Z(n483) );
  XNOR2_X1 U431 ( .A(G116), .B(G107), .ZN(n482) );
  XNOR2_X1 U432 ( .A(G143), .B(G113), .ZN(n463) );
  XNOR2_X1 U433 ( .A(G131), .B(G140), .ZN(n469) );
  INV_X1 U434 ( .A(KEYINPUT81), .ZN(n380) );
  XNOR2_X1 U435 ( .A(G902), .B(KEYINPUT15), .ZN(n381) );
  INV_X1 U436 ( .A(n730), .ZN(n393) );
  XNOR2_X1 U437 ( .A(n440), .B(n409), .ZN(n703) );
  XNOR2_X1 U438 ( .A(KEYINPUT16), .B(G122), .ZN(n409) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n702) );
  XNOR2_X1 U440 ( .A(KEYINPUT82), .B(G110), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n384), .B(G107), .ZN(n383) );
  INV_X1 U442 ( .A(G104), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n401), .B(n400), .ZN(n551) );
  XNOR2_X1 U444 ( .A(KEYINPUT28), .B(KEYINPUT103), .ZN(n400) );
  NAND2_X1 U445 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U446 ( .A(n502), .B(KEYINPUT89), .ZN(n661) );
  XNOR2_X1 U447 ( .A(n542), .B(n361), .ZN(n360) );
  XNOR2_X1 U448 ( .A(n420), .B(n365), .ZN(n699) );
  XNOR2_X1 U449 ( .A(n419), .B(n366), .ZN(n365) );
  AND2_X1 U450 ( .A1(n479), .A2(G221), .ZN(n366) );
  NAND2_X1 U451 ( .A1(n697), .A2(G478), .ZN(n604) );
  NAND2_X1 U452 ( .A1(n697), .A2(G475), .ZN(n364) );
  AND2_X2 U453 ( .A1(n616), .A2(n615), .ZN(n697) );
  XNOR2_X1 U454 ( .A(n494), .B(n359), .ZN(n495) );
  XNOR2_X1 U455 ( .A(n493), .B(n354), .ZN(n359) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n736) );
  INV_X1 U457 ( .A(KEYINPUT32), .ZN(n390) );
  NAND2_X1 U458 ( .A1(n523), .A2(n392), .ZN(n391) );
  NOR2_X1 U459 ( .A1(n590), .A2(n549), .ZN(n392) );
  AND2_X1 U460 ( .A1(n506), .A2(n657), .ZN(n627) );
  NOR2_X1 U461 ( .A1(n540), .A2(n513), .ZN(n505) );
  XNOR2_X1 U462 ( .A(n405), .B(KEYINPUT97), .ZN(n738) );
  NOR2_X1 U463 ( .A1(n407), .A2(n653), .ZN(n406) );
  INV_X1 U464 ( .A(KEYINPUT56), .ZN(n377) );
  NAND2_X1 U465 ( .A1(n379), .A2(n691), .ZN(n378) );
  XNOR2_X1 U466 ( .A(n413), .B(n614), .ZN(n379) );
  NOR2_X1 U467 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U468 ( .A1(n563), .A2(n562), .ZN(n352) );
  AND2_X1 U469 ( .A1(n394), .A2(n393), .ZN(n353) );
  AND2_X1 U470 ( .A1(G227), .A2(n726), .ZN(n354) );
  XOR2_X1 U471 ( .A(KEYINPUT22), .B(KEYINPUT65), .Z(n355) );
  XNOR2_X1 U472 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n356) );
  INV_X1 U473 ( .A(n597), .ZN(n596) );
  INV_X1 U474 ( .A(n703), .ZN(n389) );
  NAND2_X1 U475 ( .A1(n503), .A2(n492), .ZN(n357) );
  NAND2_X1 U476 ( .A1(n358), .A2(n556), .ZN(n517) );
  XNOR2_X1 U477 ( .A(n514), .B(KEYINPUT34), .ZN(n358) );
  XNOR2_X2 U478 ( .A(KEYINPUT1), .B(n550), .ZN(n649) );
  NOR2_X1 U479 ( .A1(n627), .A2(n375), .ZN(n368) );
  NAND2_X1 U480 ( .A1(n372), .A2(n371), .ZN(n370) );
  NOR2_X1 U481 ( .A1(n733), .A2(n732), .ZN(n585) );
  NAND2_X1 U482 ( .A1(n360), .A2(n543), .ZN(n544) );
  XNOR2_X1 U483 ( .A(n362), .B(n611), .ZN(G60) );
  NAND2_X1 U484 ( .A1(n363), .A2(n691), .ZN(n362) );
  XNOR2_X1 U485 ( .A(n364), .B(n610), .ZN(n363) );
  INV_X1 U486 ( .A(n653), .ZN(n549) );
  NAND2_X1 U487 ( .A1(n369), .A2(n368), .ZN(n372) );
  INV_X1 U488 ( .A(n643), .ZN(n369) );
  XNOR2_X2 U489 ( .A(n504), .B(KEYINPUT31), .ZN(n643) );
  NAND2_X1 U490 ( .A1(n643), .A2(n375), .ZN(n371) );
  NAND2_X1 U491 ( .A1(n627), .A2(n375), .ZN(n374) );
  NOR2_X1 U492 ( .A1(n682), .A2(n376), .ZN(n683) );
  NOR2_X1 U493 ( .A1(n673), .A2(n376), .ZN(n674) );
  XNOR2_X1 U494 ( .A(n378), .B(n377), .ZN(G51) );
  NOR2_X2 U495 ( .A1(n711), .A2(n724), .ZN(n686) );
  NAND2_X1 U496 ( .A1(n386), .A2(n385), .ZN(n601) );
  INV_X1 U497 ( .A(n711), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n686), .A2(KEYINPUT2), .ZN(n615) );
  XNOR2_X2 U499 ( .A(n387), .B(n450), .ZN(n571) );
  NOR2_X2 U500 ( .A1(n612), .A2(n596), .ZN(n387) );
  XNOR2_X1 U501 ( .A(n388), .B(n496), .ZN(n612) );
  XNOR2_X1 U502 ( .A(n447), .B(n389), .ZN(n388) );
  XNOR2_X2 U503 ( .A(n532), .B(n531), .ZN(n711) );
  XNOR2_X1 U504 ( .A(n505), .B(KEYINPUT86), .ZN(n506) );
  XNOR2_X2 U505 ( .A(n351), .B(n478), .ZN(n721) );
  XNOR2_X2 U506 ( .A(n721), .B(n430), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n395), .B(n588), .ZN(n394) );
  XNOR2_X2 U508 ( .A(n404), .B(n459), .ZN(n503) );
  NAND2_X1 U509 ( .A1(n408), .A2(n406), .ZN(n405) );
  XNOR2_X1 U510 ( .A(n523), .B(KEYINPUT76), .ZN(n408) );
  XNOR2_X1 U511 ( .A(n608), .B(n607), .ZN(G63) );
  XNOR2_X1 U512 ( .A(n604), .B(n603), .ZN(n606) );
  OR2_X1 U513 ( .A1(n527), .A2(n526), .ZN(n414) );
  XNOR2_X1 U514 ( .A(n441), .B(KEYINPUT18), .ZN(n443) );
  XNOR2_X1 U515 ( .A(n443), .B(n442), .ZN(n444) );
  INV_X1 U516 ( .A(n500), .ZN(n491) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT78), .ZN(n459) );
  AND2_X1 U518 ( .A1(n579), .A2(n491), .ZN(n492) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n588) );
  INV_X1 U520 ( .A(G101), .ZN(n430) );
  XNOR2_X1 U521 ( .A(KEYINPUT99), .B(KEYINPUT33), .ZN(n511) );
  INV_X1 U522 ( .A(KEYINPUT70), .ZN(n497) );
  XNOR2_X1 U523 ( .A(n497), .B(G469), .ZN(n498) );
  XNOR2_X1 U524 ( .A(n619), .B(n618), .ZN(n620) );
  INV_X1 U525 ( .A(KEYINPUT63), .ZN(n623) );
  INV_X1 U526 ( .A(n571), .ZN(n593) );
  XNOR2_X1 U527 ( .A(n623), .B(KEYINPUT109), .ZN(n624) );
  INV_X1 U528 ( .A(KEYINPUT122), .ZN(n607) );
  XNOR2_X1 U529 ( .A(n625), .B(n624), .ZN(G57) );
  XNOR2_X1 U530 ( .A(n717), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U531 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U532 ( .A(n417), .B(KEYINPUT83), .Z(n419) );
  NAND2_X1 U533 ( .A1(G234), .A2(n726), .ZN(n418) );
  NOR2_X1 U534 ( .A1(n699), .A2(G902), .ZN(n425) );
  XOR2_X1 U535 ( .A(KEYINPUT84), .B(KEYINPUT25), .Z(n423) );
  NAND2_X1 U536 ( .A1(G234), .A2(n597), .ZN(n421) );
  XNOR2_X1 U537 ( .A(KEYINPUT20), .B(n421), .ZN(n489) );
  NAND2_X1 U538 ( .A1(n489), .A2(G217), .ZN(n422) );
  XNOR2_X1 U539 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U540 ( .A(G128), .ZN(n426) );
  NAND2_X1 U541 ( .A1(G143), .A2(n426), .ZN(n429) );
  INV_X1 U542 ( .A(G143), .ZN(n427) );
  NAND2_X1 U543 ( .A1(n427), .A2(G128), .ZN(n428) );
  XNOR2_X1 U544 ( .A(G146), .B(n718), .ZN(n494) );
  XOR2_X1 U545 ( .A(n448), .B(n494), .Z(n438) );
  XNOR2_X1 U546 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U547 ( .A(n440), .B(n434), .Z(n436) );
  NOR2_X1 U548 ( .A1(G953), .A2(G237), .ZN(n460) );
  NAND2_X1 U549 ( .A1(n460), .A2(G210), .ZN(n435) );
  XNOR2_X1 U550 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U551 ( .A(n438), .B(n437), .ZN(n619) );
  NOR2_X1 U552 ( .A1(G902), .A2(n619), .ZN(n439) );
  XNOR2_X1 U553 ( .A(KEYINPUT6), .B(n657), .ZN(n570) );
  INV_X1 U554 ( .A(n444), .ZN(n446) );
  NAND2_X1 U555 ( .A1(G224), .A2(n726), .ZN(n445) );
  XNOR2_X1 U556 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U557 ( .A(KEYINPUT71), .B(n702), .ZN(n449) );
  NAND2_X1 U558 ( .A1(G210), .A2(n451), .ZN(n450) );
  NAND2_X1 U559 ( .A1(G214), .A2(n451), .ZN(n664) );
  NAND2_X1 U560 ( .A1(n571), .A2(n664), .ZN(n452) );
  NAND2_X1 U561 ( .A1(G234), .A2(G237), .ZN(n453) );
  XOR2_X1 U562 ( .A(KEYINPUT14), .B(n453), .Z(n534) );
  NAND2_X1 U563 ( .A1(G952), .A2(n726), .ZN(n533) );
  INV_X1 U564 ( .A(n533), .ZN(n455) );
  NOR2_X1 U565 ( .A1(G898), .A2(n535), .ZN(n454) );
  NOR2_X1 U566 ( .A1(n455), .A2(n454), .ZN(n456) );
  NOR2_X1 U567 ( .A1(n534), .A2(n456), .ZN(n457) );
  XNOR2_X1 U568 ( .A(KEYINPUT0), .B(KEYINPUT67), .ZN(n458) );
  NAND2_X1 U569 ( .A1(G214), .A2(n460), .ZN(n462) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n464), .B(n463), .ZN(n468) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U574 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n470) );
  XNOR2_X1 U575 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U576 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n609) );
  NOR2_X1 U578 ( .A1(G902), .A2(n609), .ZN(n476) );
  XNOR2_X1 U579 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U581 ( .A(G475), .B(n477), .Z(n516) );
  XOR2_X1 U582 ( .A(G134), .B(n478), .Z(n481) );
  NAND2_X1 U583 ( .A1(G217), .A2(n479), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n481), .B(n480), .ZN(n485) );
  XNOR2_X1 U585 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U586 ( .A(n485), .B(n484), .Z(n487) );
  XNOR2_X1 U587 ( .A(KEYINPUT96), .B(KEYINPUT7), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n602) );
  NOR2_X1 U589 ( .A1(G902), .A2(n602), .ZN(n488) );
  XOR2_X1 U590 ( .A(G478), .B(n488), .Z(n515) );
  NOR2_X1 U591 ( .A1(n516), .A2(n515), .ZN(n579) );
  NAND2_X1 U592 ( .A1(n489), .A2(G221), .ZN(n490) );
  XNOR2_X1 U593 ( .A(KEYINPUT21), .B(n490), .ZN(n654) );
  XOR2_X1 U594 ( .A(n654), .B(KEYINPUT85), .Z(n500) );
  XNOR2_X1 U595 ( .A(n496), .B(n495), .ZN(n693) );
  XNOR2_X2 U596 ( .A(n499), .B(n498), .ZN(n550) );
  INV_X1 U597 ( .A(n649), .ZN(n590) );
  NAND2_X1 U598 ( .A1(n650), .A2(n649), .ZN(n501) );
  XNOR2_X2 U599 ( .A(n501), .B(KEYINPUT73), .ZN(n510) );
  INV_X1 U600 ( .A(n657), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n510), .A2(n541), .ZN(n502) );
  NAND2_X1 U602 ( .A1(n661), .A2(n503), .ZN(n504) );
  NAND2_X1 U603 ( .A1(n550), .A2(n650), .ZN(n540) );
  INV_X1 U604 ( .A(n503), .ZN(n513) );
  INV_X1 U605 ( .A(n515), .ZN(n507) );
  AND2_X1 U606 ( .A1(n507), .A2(n516), .ZN(n639) );
  NOR2_X1 U607 ( .A1(n516), .A2(n507), .ZN(n642) );
  NOR2_X1 U608 ( .A1(n639), .A2(n642), .ZN(n670) );
  XNOR2_X1 U609 ( .A(n509), .B(KEYINPUT98), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n510), .A2(n570), .ZN(n512) );
  AND2_X1 U611 ( .A1(n516), .A2(n515), .ZN(n556) );
  XNOR2_X2 U612 ( .A(n517), .B(KEYINPUT35), .ZN(n731) );
  NAND2_X1 U613 ( .A1(n731), .A2(KEYINPUT44), .ZN(n518) );
  AND2_X1 U614 ( .A1(n519), .A2(n518), .ZN(n530) );
  NOR2_X1 U615 ( .A1(n731), .A2(KEYINPUT44), .ZN(n524) );
  NOR2_X1 U616 ( .A1(n549), .A2(n520), .ZN(n521) );
  NAND2_X1 U617 ( .A1(n521), .A2(n657), .ZN(n522) );
  NOR2_X1 U618 ( .A1(n649), .A2(n522), .ZN(n631) );
  NOR2_X1 U619 ( .A1(n631), .A2(n736), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n524), .A2(n527), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n525), .B(KEYINPUT72), .ZN(n528) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n526) );
  INV_X1 U623 ( .A(KEYINPUT45), .ZN(n531) );
  NOR2_X1 U624 ( .A1(n533), .A2(n534), .ZN(n539) );
  INV_X1 U625 ( .A(n534), .ZN(n678) );
  NOR2_X1 U626 ( .A1(G900), .A2(n535), .ZN(n536) );
  NAND2_X1 U627 ( .A1(n678), .A2(n536), .ZN(n537) );
  XOR2_X1 U628 ( .A(KEYINPUT100), .B(n537), .Z(n538) );
  NOR2_X1 U629 ( .A1(n539), .A2(n538), .ZN(n547) );
  INV_X1 U630 ( .A(n540), .ZN(n543) );
  NAND2_X1 U631 ( .A1(n541), .A2(n664), .ZN(n542) );
  NOR2_X1 U632 ( .A1(n547), .A2(n544), .ZN(n557) );
  XNOR2_X2 U633 ( .A(KEYINPUT38), .B(n593), .ZN(n665) );
  NAND2_X1 U634 ( .A1(n557), .A2(n665), .ZN(n545) );
  NAND2_X1 U635 ( .A1(n642), .A2(n576), .ZN(n546) );
  XNOR2_X1 U636 ( .A(n546), .B(KEYINPUT107), .ZN(n730) );
  NOR2_X1 U637 ( .A1(n654), .A2(n547), .ZN(n548) );
  XOR2_X1 U638 ( .A(KEYINPUT69), .B(n548), .Z(n566) );
  NAND2_X1 U639 ( .A1(n551), .A2(n550), .ZN(n582) );
  INV_X1 U640 ( .A(n582), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n553), .A2(n552), .ZN(n564) );
  NAND2_X1 U642 ( .A1(KEYINPUT74), .A2(n564), .ZN(n554) );
  INV_X1 U643 ( .A(n670), .ZN(n559) );
  NAND2_X1 U644 ( .A1(n554), .A2(n559), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n555), .A2(KEYINPUT47), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U647 ( .A1(n593), .A2(n558), .ZN(n636) );
  INV_X1 U648 ( .A(n564), .ZN(n637) );
  NAND2_X1 U649 ( .A1(n637), .A2(n559), .ZN(n560) );
  NOR2_X1 U650 ( .A1(KEYINPUT47), .A2(n560), .ZN(n561) );
  NOR2_X1 U651 ( .A1(n636), .A2(n561), .ZN(n562) );
  AND2_X1 U652 ( .A1(n564), .A2(KEYINPUT47), .ZN(n565) );
  NOR2_X1 U653 ( .A1(KEYINPUT74), .A2(n565), .ZN(n575) );
  XOR2_X1 U654 ( .A(KEYINPUT36), .B(KEYINPUT77), .Z(n573) );
  NAND2_X1 U655 ( .A1(n664), .A2(n653), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n639), .A2(n566), .ZN(n567) );
  NOR2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U658 ( .A1(n570), .A2(n569), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n589), .A2(n571), .ZN(n572) );
  XNOR2_X1 U660 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X1 U661 ( .A1(n574), .A2(n590), .ZN(n646) );
  NOR2_X1 U662 ( .A1(n575), .A2(n646), .ZN(n587) );
  XOR2_X1 U663 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n578) );
  NAND2_X1 U664 ( .A1(n576), .A2(n639), .ZN(n577) );
  XNOR2_X1 U665 ( .A(n578), .B(n577), .ZN(n733) );
  INV_X1 U666 ( .A(n579), .ZN(n667) );
  NAND2_X1 U667 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U668 ( .A1(n667), .A2(n669), .ZN(n581) );
  XOR2_X1 U669 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n580) );
  XNOR2_X1 U670 ( .A(n581), .B(n580), .ZN(n682) );
  NOR2_X1 U671 ( .A1(n682), .A2(n582), .ZN(n583) );
  XNOR2_X1 U672 ( .A(n583), .B(KEYINPUT42), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n584), .B(KEYINPUT106), .ZN(n732) );
  XNOR2_X1 U674 ( .A(n585), .B(n356), .ZN(n586) );
  XOR2_X1 U675 ( .A(n589), .B(KEYINPUT101), .Z(n591) );
  NAND2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U677 ( .A(n592), .B(KEYINPUT43), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U679 ( .A(KEYINPUT102), .B(n595), .ZN(n737) );
  NAND2_X1 U680 ( .A1(n353), .A2(n737), .ZN(n724) );
  XNOR2_X1 U681 ( .A(KEYINPUT75), .B(n597), .ZN(n598) );
  NAND2_X1 U682 ( .A1(n598), .A2(KEYINPUT2), .ZN(n599) );
  XNOR2_X1 U683 ( .A(KEYINPUT66), .B(n599), .ZN(n600) );
  XNOR2_X1 U684 ( .A(n602), .B(KEYINPUT121), .ZN(n603) );
  NOR2_X1 U685 ( .A1(G952), .A2(n726), .ZN(n605) );
  XOR2_X1 U686 ( .A(KEYINPUT80), .B(n605), .Z(n691) );
  NAND2_X1 U687 ( .A1(n606), .A2(n691), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT59), .ZN(n610) );
  INV_X1 U689 ( .A(KEYINPUT60), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT54), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT55), .ZN(n614) );
  AND2_X1 U692 ( .A1(n615), .A2(G472), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT62), .B(KEYINPUT108), .Z(n618) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n622), .A2(n691), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n627), .A2(n639), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(G104), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U700 ( .A1(n627), .A2(n642), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U702 ( .A(G107), .B(n630), .ZN(G9) );
  XNOR2_X1 U703 ( .A(G110), .B(n631), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT111), .ZN(G12) );
  XOR2_X1 U705 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n634) );
  NAND2_X1 U706 ( .A1(n637), .A2(n642), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U708 ( .A(G128), .B(n635), .ZN(G30) );
  XOR2_X1 U709 ( .A(G143), .B(n636), .Z(G45) );
  NAND2_X1 U710 ( .A1(n637), .A2(n639), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n638), .B(G146), .ZN(G48) );
  XOR2_X1 U712 ( .A(G113), .B(KEYINPUT113), .Z(n641) );
  NAND2_X1 U713 ( .A1(n643), .A2(n639), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G15) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(KEYINPUT114), .ZN(n645) );
  XNOR2_X1 U717 ( .A(G116), .B(n645), .ZN(G18) );
  XOR2_X1 U718 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n648) );
  XNOR2_X1 U719 ( .A(G125), .B(n646), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(G27) );
  XNOR2_X1 U721 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n677) );
  XOR2_X1 U722 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n652) );
  OR2_X1 U723 ( .A1(n650), .A2(n407), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT49), .B(n655), .Z(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT51), .B(n662), .Z(n663) );
  NOR2_X1 U731 ( .A1(n682), .A2(n663), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U734 ( .A(KEYINPUT117), .B(n668), .Z(n672) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U738 ( .A(n677), .B(n676), .ZN(n680) );
  NAND2_X1 U739 ( .A1(G952), .A2(n678), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U741 ( .A1(G953), .A2(n681), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n683), .B(KEYINPUT119), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n688) );
  XOR2_X1 U744 ( .A(n686), .B(KEYINPUT2), .Z(n687) );
  XNOR2_X1 U745 ( .A(n689), .B(KEYINPUT53), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n690), .B(KEYINPUT120), .ZN(G75) );
  INV_X1 U747 ( .A(n691), .ZN(n701) );
  NAND2_X1 U748 ( .A1(n697), .A2(G469), .ZN(n695) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n701), .A2(n696), .ZN(G54) );
  NAND2_X1 U753 ( .A1(G217), .A2(n697), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n701), .A2(n700), .ZN(G66) );
  XNOR2_X1 U756 ( .A(G101), .B(n702), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n706) );
  NOR2_X1 U758 ( .A1(G898), .A2(n726), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(n715) );
  INV_X1 U760 ( .A(G898), .ZN(n710) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT123), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n708), .B(KEYINPUT61), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U765 ( .A1(G953), .A2(n711), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U767 ( .A(n715), .B(n714), .Z(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT124), .B(n716), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n717), .B(KEYINPUT125), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(n725) );
  XNOR2_X1 U772 ( .A(G227), .B(n725), .ZN(n722) );
  NAND2_X1 U773 ( .A1(G900), .A2(n722), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n723), .A2(G953), .ZN(n729) );
  XNOR2_X1 U775 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U778 ( .A(G134), .B(n730), .Z(G36) );
  XOR2_X1 U779 ( .A(n731), .B(G122), .Z(G24) );
  XOR2_X1 U780 ( .A(G137), .B(n732), .Z(G39) );
  XNOR2_X1 U781 ( .A(G131), .B(n733), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U783 ( .A(G119), .B(KEYINPUT126), .Z(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(G21) );
  XNOR2_X1 U785 ( .A(G140), .B(n737), .ZN(G42) );
  XOR2_X1 U786 ( .A(n738), .B(G101), .Z(n739) );
  XNOR2_X1 U787 ( .A(KEYINPUT110), .B(n739), .ZN(G3) );
endmodule

