//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G325));
  XNOR2_X1  g033(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g034(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n465), .B1(new_n467), .B2(G101), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n462), .A2(new_n463), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n461), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n461), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n479), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n490), .B2(G114), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT72), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n462), .B2(new_n463), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n463), .C2(new_n462), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(G50), .A3(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(new_n508), .B2(new_n509), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n506), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(G89), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n504), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n522), .B(new_n523), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n528), .A2(new_n538), .B1(new_n516), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n536), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n528), .A2(new_n544), .B1(new_n516), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n510), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(G651), .A2(new_n557), .B1(new_n517), .B2(G91), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  OR2_X1    g135(.A1(new_n532), .A2(new_n533), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n505), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n563), .A2(new_n513), .A3(new_n518), .ZN(G303));
  INV_X1    g139(.A(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n524), .A2(new_n565), .A3(new_n525), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n517), .A2(G87), .B1(G651), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G49), .B(G543), .C1(new_n515), .C2(new_n514), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n504), .A2(new_n570), .A3(G49), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n567), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n579), .A2(G73), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G61), .B1(new_n508), .B2(new_n509), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n536), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n526), .A2(new_n504), .A3(G86), .ZN(new_n585));
  OAI211_X1 g160(.A(G48), .B(G543), .C1(new_n515), .C2(new_n514), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n536), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n528), .A2(new_n592), .B1(new_n516), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n510), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n515), .A2(new_n514), .ZN(new_n600));
  INV_X1    g175(.A(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n599), .A2(G651), .B1(new_n602), .B2(G54), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n516), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n516), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G171), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G171), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n609), .ZN(G280));
  XOR2_X1   g189(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g190(.A(new_n608), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n547), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n609), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n608), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g198(.A(KEYINPUT3), .B(G2104), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n467), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n461), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(KEYINPUT17), .B1(new_n653), .B2(new_n654), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n667), .A2(new_n672), .A3(new_n670), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n672), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n675));
  AOI211_X1 g250(.A(new_n671), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n674), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT83), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n681), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n679), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n688), .ZN(G229));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n588), .A2(G16), .ZN(new_n691));
  OR2_X1    g266(.A1(G6), .A2(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT32), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1981), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT84), .Z(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1971), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G23), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n567), .A2(new_n572), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n698), .A2(new_n709), .A3(KEYINPUT85), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n690), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n712), .A2(KEYINPUT86), .A3(KEYINPUT34), .A4(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n477), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n482), .A2(G119), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n461), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n699), .A2(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n595), .B2(new_n699), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n727), .B(new_n730), .C1(new_n714), .C2(new_n715), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n718), .A2(new_n731), .A3(KEYINPUT87), .A4(KEYINPUT36), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n718), .B2(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n699), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n699), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT91), .B(G1966), .Z(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G33), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n743));
  NAND2_X1  g318(.A1(G103), .A2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n477), .A2(G139), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n476), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2105), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(new_n741), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT89), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2072), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n741), .B1(KEYINPUT24), .B2(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(KEYINPUT24), .B2(G34), .ZN(new_n757));
  INV_X1    g332(.A(G160), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G27), .A2(G29), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G164), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n740), .A2(new_n755), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT90), .B1(G29), .B2(G32), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n467), .A2(G105), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n482), .A2(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n768), .B(new_n772), .C1(G141), .C2(new_n477), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  MUX2_X1   g349(.A(KEYINPUT90), .B(new_n767), .S(new_n774), .Z(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n699), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n699), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1961), .Z(new_n781));
  XOR2_X1   g356(.A(KEYINPUT31), .B(G11), .Z(new_n782));
  NOR2_X1   g357(.A1(new_n635), .A2(new_n741), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n782), .B(new_n783), .C1(new_n741), .C2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n760), .C2(new_n759), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n777), .A2(new_n778), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n737), .A2(new_n739), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT92), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n766), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT93), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n766), .A2(new_n787), .A3(new_n792), .A4(new_n789), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n741), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n741), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT29), .Z(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G4), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n616), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT88), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1348), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n699), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n547), .B2(new_n699), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n741), .A2(G26), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT28), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n477), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n482), .A2(G128), .ZN(new_n809));
  OR2_X1    g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2067), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n699), .A2(G20), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT23), .Z(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G299), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT94), .B(G1956), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n805), .B(new_n819), .C1(new_n817), .C2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n802), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n796), .B2(new_n797), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n791), .A2(new_n793), .A3(new_n798), .A4(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n733), .A2(new_n735), .A3(new_n823), .ZN(G311));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n735), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n732), .ZN(G150));
  NAND2_X1  g401(.A1(new_n616), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n510), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n536), .B1(new_n833), .B2(KEYINPUT95), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(KEYINPUT95), .B2(new_n833), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT96), .B(G55), .Z(new_n836));
  AOI22_X1  g411(.A1(G93), .A2(new_n517), .B1(new_n602), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n619), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n830), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(G860), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n838), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n846), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT99), .ZN(G145));
  XNOR2_X1  g427(.A(KEYINPUT103), .B(G37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n482), .A2(G130), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n477), .B2(G142), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n626), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n773), .B(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G164), .B(new_n812), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n723), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n635), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(G162), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n870), .A3(new_n867), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n872), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n853), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g454(.A(new_n839), .B(new_n621), .ZN(new_n880));
  OR2_X1    g455(.A1(G299), .A2(new_n608), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n608), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT104), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(KEYINPUT104), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n884), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n896));
  XNOR2_X1  g471(.A(G166), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(new_n705), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n897), .B(new_n898), .Z(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT42), .Z(new_n900));
  AND3_X1   g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g479(.A(new_n903), .B1(G868), .B2(new_n848), .ZN(G331));
  NAND2_X1  g480(.A1(G286), .A2(G301), .ZN(new_n906));
  NAND2_X1  g481(.A1(G168), .A2(G171), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n839), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n908), .B2(new_n839), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n908), .B2(new_n839), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n908), .A2(new_n839), .A3(KEYINPUT106), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n911), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n891), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n908), .A2(new_n839), .ZN(new_n917));
  OR3_X1    g492(.A1(new_n917), .A2(new_n909), .A3(new_n883), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n899), .ZN(new_n920));
  INV_X1    g495(.A(new_n899), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT43), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n917), .A2(new_n909), .B1(new_n887), .B2(new_n888), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n915), .B2(new_n883), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n899), .ZN(new_n926));
  AND4_X1   g501(.A1(KEYINPUT43), .A2(new_n926), .A3(new_n922), .A4(new_n853), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n920), .B2(new_n922), .ZN(new_n930));
  AND4_X1   g505(.A1(new_n929), .A2(new_n926), .A3(new_n922), .A4(new_n853), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n928), .B1(new_n932), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n500), .A2(new_n502), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n490), .A2(G114), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n492), .A2(KEYINPUT72), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(G2105), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n482), .A2(G126), .B1(new_n938), .B2(new_n489), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n471), .A2(new_n474), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT109), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n812), .B(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n773), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n946), .A2(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n773), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n723), .B(new_n726), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n947), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n595), .B(G1986), .Z(new_n958));
  NAND3_X1  g533(.A1(new_n943), .A2(new_n945), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n940), .A2(new_n945), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G8), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n964), .A3(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n705), .A2(G1976), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n964), .B1(new_n961), .B2(G8), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT112), .B(new_n972), .C1(new_n940), .C2(new_n945), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT52), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT49), .B1(new_n584), .B2(new_n587), .ZN(new_n976));
  INV_X1    g551(.A(G1981), .ZN(new_n977));
  INV_X1    g552(.A(G61), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n524), .B2(new_n525), .ZN(new_n979));
  OAI21_X1  g554(.A(G651), .B1(new_n979), .B2(new_n581), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n980), .B2(KEYINPUT113), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n980), .A2(new_n982), .A3(new_n585), .A4(new_n586), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n976), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n976), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n973), .B2(new_n971), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n970), .A2(new_n975), .A3(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT55), .B(G8), .C1(new_n506), .C2(new_n519), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(G166), .B2(new_n972), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  NAND4_X1  g568(.A1(G303), .A2(new_n993), .A3(KEYINPUT55), .A4(G8), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n945), .A2(new_n797), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n940), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(KEYINPUT110), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n502), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n501), .B1(new_n624), .B2(new_n498), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n495), .B(new_n494), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n471), .ZN(new_n1009));
  INV_X1    g584(.A(new_n474), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(G40), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1005), .B2(new_n934), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1971), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(G8), .B(new_n995), .C1(new_n1008), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n966), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n987), .B2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n988), .A2(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(new_n575), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n573), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(G1976), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n987), .B1(new_n974), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n966), .B2(new_n969), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1011), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT115), .B(new_n945), .C1(new_n940), .C2(new_n998), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n797), .A3(new_n999), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1013), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n945), .B1(new_n940), .B2(KEYINPUT45), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n995), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1029), .A2(new_n1042), .A3(new_n1015), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1011), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .A3(new_n760), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n738), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(G2084), .B(new_n1011), .C1(new_n1000), .C2(new_n1007), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(G168), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1022), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G168), .A2(G8), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1049), .A2(KEYINPUT116), .B1(new_n738), .B2(new_n1046), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n760), .A3(new_n945), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1015), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n988), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT117), .A4(new_n1042), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1052), .A2(new_n1053), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1053), .B1(new_n1065), .B2(new_n1041), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1060), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1021), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1033), .A2(new_n999), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n997), .B2(new_n945), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n558), .B2(KEYINPUT118), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n554), .A2(new_n1076), .A3(new_n558), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n554), .B2(new_n558), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n554), .A2(new_n1076), .A3(new_n558), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1073), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n940), .A2(new_n945), .A3(new_n948), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1044), .B2(G1348), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(new_n616), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1083), .B1(new_n1073), .B2(new_n1086), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1069), .B(new_n1087), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n616), .B2(new_n1089), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1073), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1094), .B2(new_n1091), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT60), .B(new_n1088), .C1(new_n1044), .C2(G1348), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n616), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1073), .A2(new_n1086), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1083), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .A3(new_n1087), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1097), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n1046), .B2(G1996), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1084), .A2(new_n1108), .A3(new_n950), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n961), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n547), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1100), .A2(new_n616), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1092), .B(new_n1095), .C1(new_n1106), .C2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1059), .A2(G168), .A3(new_n1047), .A4(new_n1045), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(G168), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT51), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1124), .A3(G8), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1044), .A2(KEYINPUT123), .A3(G1961), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n1044), .B2(G1961), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1012), .A2(new_n764), .A3(new_n1013), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n764), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1136), .B(new_n474), .C1(KEYINPUT124), .C2(new_n471), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1013), .B(new_n1137), .C1(KEYINPUT124), .C2(new_n471), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1134), .A2(new_n1135), .B1(new_n943), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1130), .A2(G171), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1084), .A2(KEYINPUT53), .A3(new_n764), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1044), .B2(G1961), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G301), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1127), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1127), .B1(new_n1144), .B2(G301), .ZN(new_n1147));
  OAI21_X1  g722(.A(G171), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1043), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1119), .A2(new_n1126), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1068), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1123), .A2(new_n1152), .A3(new_n1125), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1043), .A2(G301), .A3(new_n1144), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n960), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n946), .A2(G1986), .A3(G290), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n957), .A2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n953), .B(KEYINPUT46), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n949), .A2(new_n773), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n947), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n723), .A2(new_n726), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n955), .A2(new_n1171), .B1(G2067), .B2(new_n812), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n947), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1158), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(G319), .ZN(new_n1178));
  NOR3_X1   g752(.A1(G401), .A2(new_n1178), .A3(G227), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n684), .A2(new_n688), .A3(new_n1179), .ZN(new_n1180));
  OAI211_X1 g754(.A(new_n878), .B(new_n1180), .C1(new_n930), .C2(new_n931), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


