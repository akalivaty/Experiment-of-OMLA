

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765;

  INV_X1 U373 ( .A(KEYINPUT46), .ZN(n351) );
  NOR2_X1 U374 ( .A1(n762), .A2(n645), .ZN(n565) );
  XNOR2_X1 U375 ( .A(n457), .B(n367), .ZN(n695) );
  NAND2_X1 U376 ( .A1(n667), .A2(n456), .ZN(n457) );
  BUF_X1 U377 ( .A(n665), .Z(n356) );
  XNOR2_X1 U378 ( .A(n452), .B(n361), .ZN(n676) );
  XNOR2_X1 U379 ( .A(n577), .B(KEYINPUT1), .ZN(n677) );
  OR2_X1 U380 ( .A1(n632), .A2(G902), .ZN(n452) );
  NAND2_X1 U381 ( .A1(n403), .A2(n400), .ZN(n577) );
  AND2_X1 U382 ( .A1(n717), .A2(n404), .ZN(n372) );
  XNOR2_X1 U383 ( .A(n355), .B(n739), .ZN(n710) );
  XNOR2_X1 U384 ( .A(n504), .B(n419), .ZN(n355) );
  XNOR2_X1 U385 ( .A(n504), .B(n488), .ZN(n548) );
  INV_X1 U386 ( .A(G953), .ZN(n752) );
  XNOR2_X2 U387 ( .A(n454), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X2 U388 ( .A1(n559), .A2(n604), .ZN(n560) );
  XNOR2_X1 U389 ( .A(n352), .B(n351), .ZN(n384) );
  NAND2_X1 U390 ( .A1(n354), .A2(n353), .ZN(n352) );
  INV_X1 U391 ( .A(n765), .ZN(n353) );
  INV_X1 U392 ( .A(n759), .ZN(n354) );
  AND2_X2 U393 ( .A1(n473), .A2(n471), .ZN(n750) );
  NAND2_X2 U394 ( .A1(n584), .A2(n357), .ZN(n427) );
  AND2_X2 U395 ( .A1(n423), .A2(n569), .ZN(n357) );
  NOR2_X2 U396 ( .A1(n588), .A2(n578), .ZN(n640) );
  XNOR2_X2 U397 ( .A(n560), .B(KEYINPUT33), .ZN(n661) );
  XNOR2_X2 U398 ( .A(n744), .B(G101), .ZN(n504) );
  XNOR2_X1 U399 ( .A(n546), .B(n399), .ZN(n398) );
  NOR2_X2 U400 ( .A1(n574), .A2(n573), .ZN(n651) );
  INV_X1 U401 ( .A(KEYINPUT104), .ZN(n557) );
  XNOR2_X1 U402 ( .A(n470), .B(n469), .ZN(n765) );
  NOR2_X1 U403 ( .A1(n410), .A2(n409), .ZN(n408) );
  AND2_X1 U404 ( .A1(n571), .A2(n366), .ZN(n645) );
  AND2_X1 U405 ( .A1(n398), .A2(n397), .ZN(n571) );
  AND2_X1 U406 ( .A1(n398), .A2(n364), .ZN(n454) );
  OR2_X1 U407 ( .A1(n576), .A2(n450), .ZN(n447) );
  OR2_X1 U408 ( .A1(n424), .A2(n676), .ZN(n589) );
  XNOR2_X1 U409 ( .A(n721), .B(n720), .ZN(n723) );
  XOR2_X1 U410 ( .A(G125), .B(G146), .Z(n502) );
  XNOR2_X1 U411 ( .A(n371), .B(n557), .ZN(n559) );
  NAND2_X1 U412 ( .A1(n677), .A2(n678), .ZN(n371) );
  XNOR2_X1 U413 ( .A(n587), .B(KEYINPUT38), .ZN(n665) );
  INV_X1 U414 ( .A(n703), .ZN(n462) );
  OR2_X1 U415 ( .A1(n735), .A2(n370), .ZN(n445) );
  NAND2_X1 U416 ( .A1(n552), .A2(n402), .ZN(n401) );
  AND2_X1 U417 ( .A1(n606), .A2(n544), .ZN(n678) );
  XNOR2_X1 U418 ( .A(G140), .B(G131), .ZN(n547) );
  INV_X1 U419 ( .A(KEYINPUT34), .ZN(n450) );
  XNOR2_X1 U420 ( .A(n506), .B(n505), .ZN(n507) );
  BUF_X1 U421 ( .A(n577), .Z(n612) );
  XNOR2_X1 U422 ( .A(n539), .B(n538), .ZN(n572) );
  XNOR2_X1 U423 ( .A(n483), .B(n362), .ZN(n395) );
  XNOR2_X1 U424 ( .A(n376), .B(n373), .ZN(n482) );
  XNOR2_X1 U425 ( .A(KEYINPUT84), .B(KEYINPUT0), .ZN(n518) );
  OR2_X1 U426 ( .A1(G902), .A2(G237), .ZN(n509) );
  XOR2_X1 U427 ( .A(G137), .B(G134), .Z(n746) );
  XNOR2_X1 U428 ( .A(G113), .B(G143), .ZN(n528) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(n502), .Z(n749) );
  INV_X1 U430 ( .A(KEYINPUT79), .ZN(n467) );
  XNOR2_X1 U431 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n487) );
  INV_X1 U432 ( .A(KEYINPUT45), .ZN(n586) );
  NAND2_X1 U433 ( .A1(G237), .A2(G234), .ZN(n513) );
  NAND2_X1 U434 ( .A1(G214), .A2(n509), .ZN(n618) );
  XNOR2_X1 U435 ( .A(n676), .B(n451), .ZN(n558) );
  XNOR2_X1 U436 ( .A(n553), .B(KEYINPUT100), .ZN(n451) );
  XNOR2_X1 U437 ( .A(n476), .B(n474), .ZN(n606) );
  XNOR2_X1 U438 ( .A(n485), .B(n475), .ZN(n474) );
  INV_X1 U439 ( .A(KEYINPUT25), .ZN(n475) );
  XNOR2_X1 U440 ( .A(n548), .B(n468), .ZN(n717) );
  XNOR2_X1 U441 ( .A(n551), .B(n745), .ZN(n468) );
  XOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n499) );
  XNOR2_X1 U443 ( .A(KEYINPUT85), .B(KEYINPUT73), .ZN(n498) );
  XNOR2_X1 U444 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U445 ( .A1(n760), .A2(n472), .ZN(n471) );
  XNOR2_X1 U446 ( .A(n380), .B(n368), .ZN(n473) );
  INV_X1 U447 ( .A(n659), .ZN(n472) );
  BUF_X2 U448 ( .A(n735), .Z(n428) );
  NAND2_X1 U449 ( .A1(n360), .A2(n386), .ZN(n623) );
  NAND2_X1 U450 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U451 ( .A(n599), .ZN(n449) );
  INV_X1 U452 ( .A(KEYINPUT22), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n432), .B(G478), .ZN(n574) );
  OR2_X1 U454 ( .A1(n725), .A2(G902), .ZN(n432) );
  INV_X1 U455 ( .A(n594), .ZN(n425) );
  BUF_X1 U456 ( .A(n676), .Z(n438) );
  XNOR2_X1 U457 ( .A(n417), .B(n497), .ZN(n739) );
  XNOR2_X1 U458 ( .A(n495), .B(n494), .ZN(n417) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n394) );
  NOR2_X1 U461 ( .A1(G952), .A2(n752), .ZN(n730) );
  OR2_X1 U462 ( .A1(n579), .A2(n358), .ZN(n411) );
  XNOR2_X1 U463 ( .A(G137), .B(G128), .ZN(n379) );
  XOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n532) );
  XOR2_X1 U465 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n529) );
  INV_X1 U466 ( .A(n763), .ZN(n464) );
  NAND2_X1 U467 ( .A1(n455), .A2(n618), .ZN(n662) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n530) );
  XNOR2_X1 U469 ( .A(G131), .B(KEYINPUT93), .ZN(n489) );
  XOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n490) );
  XNOR2_X1 U471 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X1 U472 ( .A(KEYINPUT88), .B(G140), .ZN(n377) );
  XNOR2_X1 U473 ( .A(n481), .B(n379), .ZN(n378) );
  XNOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n481) );
  XNOR2_X1 U475 ( .A(n375), .B(n374), .ZN(n373) );
  XNOR2_X1 U476 ( .A(G110), .B(G119), .ZN(n375) );
  XNOR2_X1 U477 ( .A(KEYINPUT72), .B(KEYINPUT24), .ZN(n374) );
  NAND2_X1 U478 ( .A1(n629), .A2(n467), .ZN(n466) );
  INV_X1 U479 ( .A(KEYINPUT30), .ZN(n437) );
  XNOR2_X1 U480 ( .A(n496), .B(G107), .ZN(n550) );
  XNOR2_X1 U481 ( .A(G110), .B(G104), .ZN(n496) );
  XNOR2_X1 U482 ( .A(n459), .B(n458), .ZN(n495) );
  XNOR2_X1 U483 ( .A(G119), .B(KEYINPUT3), .ZN(n458) );
  XNOR2_X1 U484 ( .A(n460), .B(G116), .ZN(n459) );
  INV_X1 U485 ( .A(G113), .ZN(n460) );
  INV_X1 U486 ( .A(G143), .ZN(n486) );
  XNOR2_X1 U487 ( .A(G122), .B(G107), .ZN(n523) );
  XNOR2_X1 U488 ( .A(n535), .B(n441), .ZN(n719) );
  XNOR2_X1 U489 ( .A(n537), .B(n536), .ZN(n441) );
  XNOR2_X1 U490 ( .A(KEYINPUT15), .B(G902), .ZN(n629) );
  NOR2_X1 U491 ( .A1(n606), .A2(n605), .ZN(n624) );
  NOR2_X1 U492 ( .A1(n558), .A2(n603), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n503), .B(n500), .ZN(n419) );
  XNOR2_X1 U494 ( .A(n630), .B(KEYINPUT80), .ZN(n631) );
  XNOR2_X1 U495 ( .A(n622), .B(n430), .ZN(n759) );
  XNOR2_X1 U496 ( .A(n621), .B(n431), .ZN(n430) );
  INV_X1 U497 ( .A(KEYINPUT108), .ZN(n431) );
  INV_X1 U498 ( .A(KEYINPUT40), .ZN(n469) );
  INV_X1 U499 ( .A(KEYINPUT35), .ZN(n405) );
  AND2_X1 U500 ( .A1(n574), .A2(n573), .ZN(n653) );
  INV_X1 U501 ( .A(KEYINPUT92), .ZN(n434) );
  NOR2_X1 U502 ( .A1(n672), .A2(n604), .ZN(n570) );
  INV_X1 U503 ( .A(KEYINPUT124), .ZN(n391) );
  XNOR2_X1 U504 ( .A(n715), .B(n422), .ZN(n718) );
  XNOR2_X1 U505 ( .A(n717), .B(n716), .ZN(n422) );
  OR2_X1 U506 ( .A1(n663), .A2(n442), .ZN(n358) );
  INV_X1 U507 ( .A(n618), .ZN(n424) );
  XNOR2_X1 U508 ( .A(KEYINPUT103), .B(n554), .ZN(n359) );
  AND2_X1 U509 ( .A1(n390), .A2(n389), .ZN(n360) );
  XOR2_X1 U510 ( .A(KEYINPUT70), .B(G472), .Z(n361) );
  NAND2_X1 U511 ( .A1(n525), .A2(G221), .ZN(n362) );
  AND2_X1 U512 ( .A1(n412), .A2(n411), .ZN(n363) );
  INV_X1 U513 ( .A(n606), .ZN(n672) );
  AND2_X1 U514 ( .A1(n555), .A2(n359), .ZN(n364) );
  AND2_X1 U515 ( .A1(n404), .A2(G902), .ZN(n365) );
  AND2_X1 U516 ( .A1(n438), .A2(n672), .ZN(n366) );
  BUF_X1 U517 ( .A(n677), .Z(n420) );
  INV_X1 U518 ( .A(n420), .ZN(n397) );
  XOR2_X1 U519 ( .A(KEYINPUT41), .B(n619), .Z(n367) );
  INV_X1 U520 ( .A(G902), .ZN(n402) );
  XOR2_X1 U521 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n368) );
  OR2_X1 U522 ( .A1(n629), .A2(n628), .ZN(n369) );
  OR2_X1 U523 ( .A1(n629), .A2(n467), .ZN(n370) );
  INV_X1 U524 ( .A(KEYINPUT102), .ZN(n442) );
  AND2_X2 U525 ( .A1(n463), .A2(n462), .ZN(n729) );
  NAND2_X1 U526 ( .A1(n729), .A2(G217), .ZN(n396) );
  NOR2_X1 U527 ( .A1(n371), .A2(n438), .ZN(n684) );
  AND2_X1 U528 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U529 ( .A1(n447), .A2(n449), .ZN(n409) );
  NOR2_X1 U530 ( .A1(n372), .A2(n365), .ZN(n403) );
  NOR2_X1 U531 ( .A1(n661), .A2(n450), .ZN(n410) );
  NAND2_X1 U532 ( .A1(n395), .A2(n402), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n384), .A2(n381), .ZN(n380) );
  NOR2_X1 U534 ( .A1(n382), .A2(n617), .ZN(n381) );
  NAND2_X1 U535 ( .A1(n383), .A2(n464), .ZN(n382) );
  INV_X1 U536 ( .A(n656), .ZN(n383) );
  NAND2_X1 U537 ( .A1(n623), .A2(n651), .ZN(n470) );
  NOR2_X1 U538 ( .A1(n356), .A2(KEYINPUT39), .ZN(n387) );
  INV_X1 U539 ( .A(n598), .ZN(n388) );
  NAND2_X1 U540 ( .A1(n665), .A2(KEYINPUT39), .ZN(n389) );
  NAND2_X1 U541 ( .A1(n598), .A2(KEYINPUT39), .ZN(n390) );
  NAND2_X1 U542 ( .A1(n595), .A2(n436), .ZN(n598) );
  XNOR2_X1 U543 ( .A(n392), .B(n391), .ZN(G66) );
  NAND2_X1 U544 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X1 U545 ( .A(n730), .ZN(n393) );
  OR2_X1 U546 ( .A1(n717), .A2(n401), .ZN(n400) );
  INV_X1 U547 ( .A(n552), .ZN(n404) );
  XNOR2_X2 U548 ( .A(n406), .B(n405), .ZN(n580) );
  NAND2_X1 U549 ( .A1(n408), .A2(n407), .ZN(n406) );
  NAND2_X1 U550 ( .A1(n448), .A2(n661), .ZN(n407) );
  NAND2_X1 U551 ( .A1(n761), .A2(KEYINPUT102), .ZN(n412) );
  XNOR2_X2 U552 ( .A(n429), .B(KEYINPUT101), .ZN(n761) );
  NAND2_X1 U553 ( .A1(n363), .A2(n413), .ZN(n416) );
  NAND2_X1 U554 ( .A1(n415), .A2(n414), .ZN(n413) );
  NOR2_X1 U555 ( .A1(n761), .A2(KEYINPUT102), .ZN(n414) );
  OR2_X1 U556 ( .A1(n579), .A2(n663), .ZN(n415) );
  NOR2_X1 U557 ( .A1(n416), .A2(n583), .ZN(n584) );
  XNOR2_X2 U558 ( .A(n519), .B(n487), .ZN(n744) );
  AND2_X1 U559 ( .A1(n443), .A2(n465), .ZN(n444) );
  BUF_X1 U560 ( .A(n587), .Z(n421) );
  NOR2_X2 U561 ( .A1(n428), .A2(n631), .ZN(n703) );
  NOR2_X1 U562 ( .A1(n580), .A2(KEYINPUT81), .ZN(n563) );
  XNOR2_X1 U563 ( .A(n510), .B(n511), .ZN(n614) );
  AND2_X1 U564 ( .A1(n750), .A2(n466), .ZN(n465) );
  NAND2_X1 U565 ( .A1(n566), .A2(n567), .ZN(n568) );
  NAND2_X1 U566 ( .A1(n576), .A2(n545), .ZN(n546) );
  NAND2_X1 U567 ( .A1(n561), .A2(n562), .ZN(n423) );
  AND2_X1 U568 ( .A1(n576), .A2(n425), .ZN(n435) );
  XNOR2_X2 U569 ( .A(n453), .B(n518), .ZN(n576) );
  NOR2_X2 U570 ( .A1(n635), .A2(n730), .ZN(n637) );
  XNOR2_X1 U571 ( .A(n426), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U572 ( .A1(n724), .A2(n730), .ZN(n426) );
  XNOR2_X2 U573 ( .A(n427), .B(n586), .ZN(n735) );
  XNOR2_X1 U574 ( .A(n482), .B(n749), .ZN(n483) );
  NAND2_X1 U575 ( .A1(n444), .A2(n445), .ZN(n461) );
  NAND2_X1 U576 ( .A1(n461), .A2(n369), .ZN(n463) );
  NAND2_X1 U577 ( .A1(n571), .A2(n570), .ZN(n429) );
  XNOR2_X1 U578 ( .A(n524), .B(n433), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n519), .B(n523), .ZN(n433) );
  XNOR2_X1 U580 ( .A(n435), .B(n434), .ZN(n578) );
  XNOR2_X1 U581 ( .A(n589), .B(n437), .ZN(n436) );
  XNOR2_X1 U582 ( .A(n439), .B(n607), .ZN(n608) );
  AND2_X1 U583 ( .A1(n421), .A2(n624), .ZN(n439) );
  NAND2_X1 U584 ( .A1(n651), .A2(n440), .ZN(n605) );
  NAND2_X1 U585 ( .A1(n735), .A2(n467), .ZN(n443) );
  XNOR2_X2 U586 ( .A(n446), .B(n486), .ZN(n519) );
  XNOR2_X2 U587 ( .A(G128), .B(KEYINPUT75), .ZN(n446) );
  AND2_X1 U588 ( .A1(n576), .A2(n450), .ZN(n448) );
  NOR2_X2 U589 ( .A1(n614), .A2(n517), .ZN(n453) );
  INV_X1 U590 ( .A(n665), .ZN(n455) );
  INV_X1 U591 ( .A(n662), .ZN(n456) );
  INV_X1 U592 ( .A(n580), .ZN(n581) );
  XNOR2_X1 U593 ( .A(n580), .B(G122), .ZN(G24) );
  NOR2_X2 U594 ( .A1(n713), .A2(n730), .ZN(n714) );
  AND2_X1 U595 ( .A1(n530), .A2(G210), .ZN(n477) );
  INV_X1 U596 ( .A(KEYINPUT65), .ZN(n564) );
  BUF_X1 U597 ( .A(n661), .Z(n693) );
  XNOR2_X1 U598 ( .A(n491), .B(n477), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n746), .B(G146), .ZN(n488) );
  INV_X1 U600 ( .A(KEYINPUT76), .ZN(n505) );
  XNOR2_X1 U601 ( .A(n492), .B(n495), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n548), .B(n493), .ZN(n632) );
  XOR2_X1 U603 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n479) );
  NAND2_X1 U604 ( .A1(G234), .A2(n752), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U606 ( .A(KEYINPUT78), .B(n480), .Z(n525) );
  NAND2_X1 U607 ( .A1(n629), .A2(G234), .ZN(n484) );
  XNOR2_X1 U608 ( .A(n484), .B(KEYINPUT20), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n540), .A2(G217), .ZN(n485) );
  XOR2_X1 U610 ( .A(n490), .B(n489), .Z(n491) );
  INV_X1 U611 ( .A(KEYINPUT19), .ZN(n511) );
  INV_X1 U612 ( .A(n550), .ZN(n497) );
  XNOR2_X1 U613 ( .A(n499), .B(n498), .ZN(n500) );
  AND2_X1 U614 ( .A1(G224), .A2(n752), .ZN(n501) );
  NAND2_X1 U615 ( .A1(n710), .A2(n629), .ZN(n508) );
  NAND2_X1 U616 ( .A1(G210), .A2(n509), .ZN(n506) );
  XNOR2_X2 U617 ( .A(n508), .B(n507), .ZN(n587) );
  NAND2_X1 U618 ( .A1(n587), .A2(n618), .ZN(n510) );
  NOR2_X1 U619 ( .A1(G898), .A2(n752), .ZN(n741) );
  NAND2_X1 U620 ( .A1(G902), .A2(n741), .ZN(n512) );
  NAND2_X1 U621 ( .A1(G952), .A2(n752), .ZN(n591) );
  NAND2_X1 U622 ( .A1(n512), .A2(n591), .ZN(n516) );
  XOR2_X1 U623 ( .A(KEYINPUT86), .B(KEYINPUT14), .Z(n514) );
  XNOR2_X1 U624 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U625 ( .A(KEYINPUT71), .B(n515), .ZN(n660) );
  NAND2_X1 U626 ( .A1(n516), .A2(n660), .ZN(n517) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n521) );
  XNOR2_X1 U628 ( .A(G116), .B(G134), .ZN(n520) );
  XNOR2_X1 U629 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U630 ( .A(n522), .B(KEYINPUT98), .Z(n524) );
  NAND2_X1 U631 ( .A1(G217), .A2(n525), .ZN(n526) );
  XNOR2_X1 U632 ( .A(n527), .B(n526), .ZN(n725) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(G475), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n534) );
  NAND2_X1 U635 ( .A1(n530), .A2(G214), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U637 ( .A(n534), .B(n533), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n547), .B(G104), .ZN(n536) );
  XNOR2_X1 U639 ( .A(n749), .B(G122), .ZN(n535) );
  NOR2_X1 U640 ( .A1(G902), .A2(n719), .ZN(n538) );
  NOR2_X1 U641 ( .A1(n574), .A2(n572), .ZN(n667) );
  XOR2_X1 U642 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n542) );
  NAND2_X1 U643 ( .A1(n540), .A2(G221), .ZN(n541) );
  XNOR2_X1 U644 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U645 ( .A(KEYINPUT90), .B(n543), .ZN(n673) );
  INV_X1 U646 ( .A(n673), .ZN(n544) );
  AND2_X1 U647 ( .A1(n667), .A2(n544), .ZN(n545) );
  XNOR2_X1 U648 ( .A(KEYINPUT87), .B(n547), .ZN(n745) );
  AND2_X1 U649 ( .A1(G227), .A2(n752), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U651 ( .A(KEYINPUT69), .B(G469), .ZN(n552) );
  INV_X1 U652 ( .A(KEYINPUT6), .ZN(n553) );
  XNOR2_X1 U653 ( .A(KEYINPUT74), .B(n558), .ZN(n555) );
  NAND2_X1 U654 ( .A1(n672), .A2(n420), .ZN(n554) );
  INV_X1 U655 ( .A(KEYINPUT44), .ZN(n556) );
  AND2_X1 U656 ( .A1(n565), .A2(n556), .ZN(n562) );
  INV_X1 U657 ( .A(n558), .ZN(n604) );
  NAND2_X1 U658 ( .A1(n574), .A2(n572), .ZN(n599) );
  XNOR2_X1 U659 ( .A(n580), .B(n564), .ZN(n561) );
  INV_X1 U660 ( .A(n563), .ZN(n567) );
  NAND2_X1 U661 ( .A1(n568), .A2(KEYINPUT44), .ZN(n569) );
  XNOR2_X1 U662 ( .A(n572), .B(KEYINPUT97), .ZN(n573) );
  XOR2_X1 U663 ( .A(KEYINPUT99), .B(n653), .Z(n596) );
  NOR2_X1 U664 ( .A1(n651), .A2(n596), .ZN(n663) );
  NAND2_X1 U665 ( .A1(n684), .A2(n576), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n575), .B(KEYINPUT31), .ZN(n654) );
  INV_X1 U667 ( .A(n438), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n612), .A2(n678), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n654), .A2(n640), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n581), .A2(KEYINPUT44), .ZN(n582) );
  AND2_X1 U671 ( .A1(n582), .A2(KEYINPUT81), .ZN(n583) );
  NOR2_X1 U672 ( .A1(G900), .A2(n752), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n590), .A2(G902), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U675 ( .A1(n593), .A2(n660), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n594), .A2(n602), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n623), .ZN(n597) );
  XNOR2_X1 U678 ( .A(KEYINPUT111), .B(n597), .ZN(n760) );
  INV_X1 U679 ( .A(n421), .ZN(n626) );
  NOR2_X1 U680 ( .A1(n599), .A2(n626), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n388), .A2(n600), .ZN(n601) );
  XNOR2_X1 U682 ( .A(KEYINPUT105), .B(n601), .ZN(n763) );
  XOR2_X1 U683 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n607) );
  NOR2_X1 U684 ( .A1(n673), .A2(n602), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n609), .A2(n618), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n397), .A2(n608), .ZN(n656) );
  NAND2_X1 U687 ( .A1(n672), .A2(n609), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n676), .A2(n610), .ZN(n611) );
  XNOR2_X1 U689 ( .A(KEYINPUT28), .B(n611), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n614), .A2(n620), .ZN(n648) );
  INV_X1 U692 ( .A(n663), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n648), .A2(n615), .ZN(n616) );
  XNOR2_X1 U694 ( .A(KEYINPUT47), .B(n616), .ZN(n617) );
  XOR2_X1 U695 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n619) );
  NOR2_X1 U696 ( .A1(n695), .A2(n620), .ZN(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n397), .A2(n624), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT43), .B(n625), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n659) );
  INV_X1 U701 ( .A(n750), .ZN(n700) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n750), .A2(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n729), .A2(G472), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT62), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT63), .B(KEYINPUT82), .Z(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(G57) );
  NAND2_X1 U709 ( .A1(n640), .A2(n651), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT112), .ZN(n639) );
  XNOR2_X1 U711 ( .A(G104), .B(n639), .ZN(G6) );
  XOR2_X1 U712 ( .A(G107), .B(KEYINPUT113), .Z(n642) );
  NAND2_X1 U713 ( .A1(n640), .A2(n653), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n644) );
  XOR2_X1 U715 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(G9) );
  XOR2_X1 U717 ( .A(G110), .B(n645), .Z(G12) );
  XOR2_X1 U718 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n653), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G30) );
  XOR2_X1 U721 ( .A(G146), .B(KEYINPUT115), .Z(n650) );
  NAND2_X1 U722 ( .A1(n648), .A2(n651), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(G48) );
  NAND2_X1 U724 ( .A1(n654), .A2(n651), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(G113), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(G116), .ZN(G18) );
  XNOR2_X1 U728 ( .A(n656), .B(KEYINPUT116), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT37), .ZN(n658) );
  XNOR2_X1 U730 ( .A(G125), .B(n658), .ZN(G27) );
  XNOR2_X1 U731 ( .A(G140), .B(n659), .ZN(G42) );
  NAND2_X1 U732 ( .A1(G952), .A2(n660), .ZN(n692) );
  NOR2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT119), .ZN(n669) );
  NAND2_X1 U735 ( .A1(n424), .A2(n356), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n693), .A2(n670), .ZN(n671) );
  XOR2_X1 U739 ( .A(KEYINPUT120), .B(n671), .Z(n689) );
  AND2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(KEYINPUT49), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n438), .A2(n675), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n678), .A2(n420), .ZN(n679) );
  XNOR2_X1 U744 ( .A(n679), .B(KEYINPUT50), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(n682), .Z(n683) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(n685), .Z(n686) );
  NOR2_X1 U749 ( .A1(n695), .A2(n686), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n687), .B(KEYINPUT118), .ZN(n688) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U754 ( .A(n693), .ZN(n694) );
  NOR2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U757 ( .A(KEYINPUT121), .B(n698), .Z(n699) );
  NAND2_X1 U758 ( .A1(n699), .A2(n752), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n428), .A2(n700), .ZN(n701) );
  NOR2_X1 U760 ( .A1(KEYINPUT2), .A2(n701), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U764 ( .A(KEYINPUT83), .B(KEYINPUT77), .Z(n708) );
  XNOR2_X1 U765 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U767 ( .A(n710), .B(n709), .Z(n712) );
  NAND2_X1 U768 ( .A1(n729), .A2(G210), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n711), .B(n712), .ZN(n713) );
  XNOR2_X1 U770 ( .A(n714), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n716) );
  NAND2_X1 U772 ( .A1(n729), .A2(G469), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n730), .A2(n718), .ZN(G54) );
  XOR2_X1 U774 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n721) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT64), .ZN(n720) );
  NAND2_X1 U776 ( .A1(n729), .A2(G475), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n722), .B(n723), .ZN(n724) );
  XOR2_X1 U778 ( .A(n725), .B(KEYINPUT123), .Z(n727) );
  NAND2_X1 U779 ( .A1(n729), .A2(G478), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n730), .A2(n728), .ZN(G63) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n732) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(G898), .A2(n733), .ZN(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT126), .B(n734), .Z(n737) );
  NOR2_X1 U787 ( .A1(G953), .A2(n428), .ZN(n736) );
  NOR2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n738), .B(KEYINPUT127), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n739), .B(G101), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(G69) );
  XOR2_X1 U793 ( .A(n746), .B(n745), .Z(n747) );
  XNOR2_X1 U794 ( .A(n744), .B(n747), .ZN(n748) );
  XNOR2_X1 U795 ( .A(n749), .B(n748), .ZN(n754) );
  INV_X1 U796 ( .A(n754), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n751), .B(n750), .ZN(n753) );
  NAND2_X1 U798 ( .A1(n753), .A2(n752), .ZN(n758) );
  XNOR2_X1 U799 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U800 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U801 ( .A1(n756), .A2(G953), .ZN(n757) );
  NAND2_X1 U802 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U803 ( .A(n759), .B(G137), .Z(G39) );
  XOR2_X1 U804 ( .A(G134), .B(n760), .Z(G36) );
  XOR2_X1 U805 ( .A(n761), .B(G101), .Z(G3) );
  XOR2_X1 U806 ( .A(n762), .B(G119), .Z(G21) );
  XOR2_X1 U807 ( .A(G143), .B(n763), .Z(n764) );
  XNOR2_X1 U808 ( .A(KEYINPUT114), .B(n764), .ZN(G45) );
  XOR2_X1 U809 ( .A(n765), .B(G131), .Z(G33) );
endmodule

