//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n215), .B1(new_n208), .B2(new_n209), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n216), .A2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G58), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  INV_X1    g0041(.A(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G1698), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n248), .A2(G223), .B1(G77), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n256), .B2(new_n257), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n262), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT67), .B(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n263), .A2(new_n264), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n259), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n267), .A2(new_n269), .B1(new_n272), .B2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n260), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G169), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n211), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n278), .A2(new_n280), .A3(G13), .A4(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n270), .A2(new_n285), .A3(G13), .A4(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n210), .B1(new_n205), .B2(new_n243), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n282), .B1(new_n290), .B2(KEYINPUT69), .ZN(new_n291));
  AOI211_X1 g0091(.A(KEYINPUT69), .B(new_n288), .C1(new_n284), .C2(new_n286), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(G50), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n287), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n297));
  INV_X1    g0097(.A(G150), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n211), .A2(new_n243), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n211), .A2(G33), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n297), .B1(new_n298), .B2(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n295), .A2(new_n296), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n274), .A2(G179), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n276), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n290), .A2(new_n308), .A3(new_n282), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n300), .A2(new_n299), .B1(new_n211), .B2(new_n308), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n288), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G77), .B2(new_n287), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n253), .A2(G232), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n248), .A2(G238), .B1(G107), .B2(new_n251), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n258), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n272), .A2(G244), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n267), .A2(new_n269), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n325), .B2(G190), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n321), .B2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR3_X1    g0128(.A1(new_n321), .A2(G179), .A3(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n321), .B2(new_n324), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n316), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n275), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT71), .B1(new_n274), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n294), .B2(new_n303), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n338), .B(new_n344), .C1(new_n339), .C2(new_n341), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n307), .B(new_n333), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  INV_X1    g0147(.A(G87), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n247), .A2(new_n347), .B1(new_n243), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G1698), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n246), .A2(G223), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n253), .A2(KEYINPUT79), .A3(G223), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT80), .B1(new_n355), .B2(new_n258), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT80), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n354), .A2(new_n353), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n259), .C1(new_n358), .C2(new_n349), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n272), .A2(G232), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n323), .A3(new_n336), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n355), .A2(new_n258), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n323), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n334), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT76), .ZN(new_n368));
  AND3_X1   g0168(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT75), .B1(G58), .B2(G68), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n211), .B1(new_n371), .B2(new_n202), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n299), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n369), .A2(new_n370), .A3(new_n201), .ZN(new_n376));
  OAI221_X1 g0176(.A(KEYINPUT76), .B1(new_n373), .B2(new_n299), .C1(new_n376), .C2(new_n211), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n251), .B2(new_n211), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n249), .A2(new_n250), .A3(new_n379), .A4(G20), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT16), .A4(new_n381), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n288), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n300), .ZN(new_n387));
  INV_X1    g0187(.A(new_n282), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n288), .B1(new_n284), .B2(new_n286), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT69), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n292), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n295), .A2(new_n387), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n392), .B2(new_n395), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n367), .B(new_n386), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT17), .ZN(new_n399));
  AOI22_X1  g0199(.A1(G238), .A2(new_n272), .B1(new_n267), .B2(new_n269), .ZN(new_n400));
  AND2_X1   g0200(.A1(G232), .A2(G1698), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n246), .A2(new_n401), .B1(G33), .B2(G97), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n350), .A2(G226), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n251), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n246), .A2(KEYINPUT72), .A3(G226), .A4(new_n350), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n259), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT73), .B1(new_n407), .B2(new_n259), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n400), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n400), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  INV_X1    g0215(.A(G68), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G20), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(new_n301), .B2(new_n308), .C1(new_n296), .C2(new_n299), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n288), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n282), .A2(new_n416), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n389), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n295), .A2(new_n416), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n411), .A2(G190), .A3(new_n413), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n415), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n407), .A2(new_n259), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n259), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n412), .B1(new_n436), .B2(new_n400), .ZN(new_n437));
  INV_X1    g0237(.A(new_n413), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n431), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT14), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n414), .A2(KEYINPUT74), .A3(new_n431), .A4(G169), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n411), .A2(G179), .A3(new_n413), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n441), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n430), .B1(new_n446), .B2(new_n426), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n386), .B1(new_n396), .B2(new_n397), .ZN(new_n448));
  INV_X1    g0248(.A(G179), .ZN(new_n449));
  INV_X1    g0249(.A(new_n365), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n356), .A2(new_n359), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n330), .B1(new_n364), .B2(new_n365), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(new_n453), .A3(KEYINPUT81), .A4(KEYINPUT18), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT18), .ZN(new_n458));
  INV_X1    g0258(.A(new_n386), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n300), .B1(new_n291), .B2(new_n293), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT78), .B1(new_n460), .B2(new_n394), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n451), .A2(new_n452), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n457), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n346), .A2(new_n399), .A3(new_n447), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n278), .A2(new_n280), .A3(G45), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G270), .B(new_n258), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n262), .A2(new_n270), .A3(new_n473), .A4(G45), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT86), .A2(G303), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT86), .A2(G303), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n244), .B(new_n245), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n350), .C1(new_n249), .C2(new_n250), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n482), .A2(new_n483), .A3(new_n259), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n482), .B2(new_n259), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n270), .A2(G33), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n287), .A2(G116), .A3(new_n289), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G33), .A3(G283), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n211), .B1(new_n494), .B2(G33), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n497), .A2(KEYINPUT20), .A3(new_n288), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n495), .B1(new_n490), .B2(new_n492), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n288), .A2(new_n499), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n284), .A2(new_n286), .A3(new_n498), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n488), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n486), .A2(new_n507), .A3(G169), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n485), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n482), .A2(new_n483), .A3(new_n259), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n475), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G179), .A3(new_n507), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n486), .A2(new_n507), .A3(KEYINPUT21), .A4(G169), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n507), .B1(G200), .B2(new_n486), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(G190), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n246), .A2(G238), .A3(new_n350), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G116), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  OAI211_X1 g0323(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n523), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n259), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G250), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n259), .B1(new_n468), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n468), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n261), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n524), .A2(new_n523), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n526), .A3(new_n522), .A4(new_n521), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n259), .B1(new_n532), .B2(new_n530), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G190), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n211), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n348), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n211), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n301), .B2(new_n494), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n288), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n284), .A2(new_n286), .A3(new_n311), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n389), .A2(G87), .A3(new_n487), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n535), .A2(new_n539), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT88), .B1(new_n522), .B2(G20), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT88), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n211), .A3(G33), .A4(G116), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(G20), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n211), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n246), .A2(new_n565), .A3(new_n211), .A4(G87), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n288), .B1(new_n567), .B2(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n569), .B(new_n562), .C1(new_n564), .C2(new_n566), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n389), .A2(G107), .A3(new_n487), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT25), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(KEYINPUT89), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n287), .B2(G107), .ZN(new_n575));
  XNOR2_X1  g0375(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n284), .A2(new_n286), .A3(new_n560), .A4(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n572), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n246), .A2(G257), .A3(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n246), .A2(G250), .A3(new_n350), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G294), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n259), .B1(new_n531), .B2(new_n473), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n259), .A2(new_n582), .B1(new_n583), .B2(G264), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(G190), .A3(new_n474), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n259), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(G264), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n474), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n571), .A2(new_n578), .A3(new_n585), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n534), .A2(new_n330), .ZN(new_n591));
  INV_X1    g0391(.A(new_n311), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n389), .A2(new_n592), .A3(new_n487), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n551), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n528), .A2(new_n449), .A3(new_n533), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n588), .A2(new_n330), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n584), .A2(new_n449), .A3(new_n474), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n568), .A2(new_n570), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n572), .A2(new_n575), .A3(new_n577), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n554), .A2(new_n590), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G244), .B(new_n350), .C1(new_n249), .C2(new_n250), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n246), .A2(KEYINPUT4), .A3(G244), .A4(new_n350), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n246), .A2(G250), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n493), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n259), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(new_n258), .C1(new_n468), .C2(new_n471), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n474), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n330), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n211), .A2(new_n243), .A3(G77), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(new_n494), .A3(G107), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n211), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n379), .B1(new_n246), .B2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n560), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n288), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n389), .A2(G97), .A3(new_n487), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n295), .A2(new_n494), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n610), .A2(new_n628), .A3(new_n474), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n610), .B2(new_n474), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n609), .B(new_n449), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n614), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n609), .A2(G190), .A3(new_n612), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n625), .A3(new_n624), .A4(new_n626), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n629), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n334), .B1(new_n637), .B2(new_n609), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT84), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n609), .B1(new_n630), .B2(new_n631), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT84), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n634), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n633), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n520), .A2(new_n602), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n467), .A2(new_n646), .ZN(G372));
  NOR3_X1   g0447(.A1(new_n463), .A2(new_n458), .A3(new_n464), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT18), .B1(new_n448), .B2(new_n453), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT92), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n465), .A2(new_n651), .A3(new_n454), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n329), .A2(new_n316), .A3(new_n331), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n446), .A2(new_n426), .B1(new_n429), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n399), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n343), .A2(new_n345), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n307), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT93), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  AOI211_X1 g0463(.A(new_n663), .B(new_n307), .C1(new_n657), .C2(new_n658), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n467), .ZN(new_n667));
  INV_X1    g0467(.A(new_n596), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n510), .A2(new_n601), .A3(new_n514), .A4(new_n515), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n551), .A2(KEYINPUT90), .A3(new_n552), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT90), .B1(new_n551), .B2(new_n552), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n535), .B(new_n539), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n596), .A3(new_n590), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n674), .B2(new_n645), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n554), .A2(new_n596), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n633), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n633), .A3(new_n596), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n633), .A2(new_n554), .A3(new_n596), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n666), .A2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(G13), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n270), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n507), .A2(new_n695), .ZN(new_n696));
  MUX2_X1   g0496(.A(new_n516), .B(new_n520), .S(new_n696), .Z(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n601), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n695), .B1(new_n599), .B2(new_n600), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n590), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n601), .A2(new_n695), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n695), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n704), .A2(new_n516), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n708), .ZN(G399));
  NAND3_X1  g0509(.A1(new_n542), .A2(new_n348), .A3(new_n498), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  INV_X1    g0511(.A(new_n206), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n711), .A2(new_n277), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n214), .B2(new_n713), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n538), .A2(new_n609), .A3(new_n612), .A4(new_n584), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n513), .A2(G179), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT95), .B(KEYINPUT30), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n718), .B2(new_n719), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n584), .B2(new_n474), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n486), .A3(new_n640), .A4(new_n534), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(KEYINPUT96), .A3(new_n725), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n717), .B(new_n706), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n721), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n717), .A3(new_n723), .A4(new_n725), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n646), .A2(KEYINPUT31), .B1(new_n732), .B2(new_n695), .ZN(new_n733));
  OAI21_X1  g0533(.A(G330), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n685), .A2(new_n706), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n639), .A2(new_n644), .ZN(new_n739));
  INV_X1    g0539(.A(new_n633), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n645), .A2(KEYINPUT97), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n674), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n596), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .A3(new_n706), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n735), .B1(new_n738), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n716), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n277), .B1(new_n689), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n713), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n699), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G330), .B2(new_n697), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n210), .B1(G20), .B2(new_n330), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n211), .A2(new_n449), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G190), .A3(new_n334), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n211), .A2(G179), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n761), .A2(G322), .B1(new_n765), .B2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n759), .A2(new_n763), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n766), .B(new_n251), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n759), .A2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n336), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(G326), .B1(new_n773), .B2(G303), .ZN(new_n774));
  INV_X1    g0574(.A(G294), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n336), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n211), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n770), .A2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT33), .B(G317), .Z(new_n780));
  OAI221_X1 g0580(.A(new_n774), .B1(new_n775), .B2(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n762), .A2(new_n336), .A3(G200), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT98), .Z(new_n783));
  AOI211_X1 g0583(.A(new_n769), .B(new_n781), .C1(G283), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n783), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n560), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n777), .A2(new_n494), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n765), .A2(G159), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(KEYINPUT32), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n251), .B1(new_n761), .B2(G58), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(new_n308), .C2(new_n768), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n778), .A2(G68), .B1(new_n773), .B2(G87), .ZN(new_n792));
  INV_X1    g0592(.A(new_n771), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(KEYINPUT32), .B2(new_n788), .C1(new_n296), .C2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n786), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n758), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n755), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n758), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n712), .A2(new_n251), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G355), .B1(new_n498), .B2(new_n712), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n237), .A2(new_n264), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n712), .A2(new_n246), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G45), .B2(new_n213), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n797), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n800), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n697), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n757), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND4_X1  g0612(.A1(new_n329), .A2(new_n316), .A3(new_n331), .A4(new_n706), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n315), .A2(new_n706), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n326), .B2(new_n327), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n654), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n736), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n682), .A2(new_n678), .A3(new_n680), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n679), .A2(new_n680), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT91), .ZN(new_n821));
  INV_X1    g0621(.A(new_n683), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n510), .A2(new_n601), .A3(new_n514), .A4(new_n515), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n824), .A2(new_n596), .A3(new_n590), .A4(new_n672), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n596), .B1(new_n825), .B2(new_n741), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n818), .B(new_n706), .C1(new_n823), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n817), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n755), .B1(new_n828), .B2(new_n734), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n735), .A2(new_n817), .A3(new_n827), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n779), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n787), .B(new_n833), .C1(G303), .C2(new_n771), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n251), .B1(new_n772), .B2(new_n560), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT99), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n783), .A2(G87), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n768), .A2(new_n498), .B1(new_n764), .B2(new_n767), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G294), .B2(new_n761), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  INV_X1    g0641(.A(G58), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n246), .B1(new_n764), .B2(new_n841), .C1(new_n777), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n785), .A2(new_n416), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(G50), .C2(new_n773), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  INV_X1    g0647(.A(new_n768), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n761), .A2(G143), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n779), .B2(new_n298), .C1(new_n850), .C2(new_n793), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT34), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n840), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n758), .ZN(new_n856));
  INV_X1    g0656(.A(new_n755), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n758), .A2(new_n798), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n308), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n798), .B2(new_n816), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n831), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NOR2_X1   g0663(.A1(new_n270), .A2(new_n689), .ZN(new_n864));
  INV_X1    g0664(.A(G330), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n646), .A2(KEYINPUT31), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n732), .A2(new_n695), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT31), .B(new_n695), .C1(new_n726), .C2(new_n721), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n667), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT107), .Z(new_n872));
  NOR2_X1   g0672(.A1(new_n396), .A2(new_n397), .ZN(new_n873));
  INV_X1    g0673(.A(new_n385), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n382), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT104), .A4(new_n381), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n383), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n288), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(KEYINPUT105), .ZN(new_n880));
  INV_X1    g0680(.A(new_n383), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n382), .B2(new_n875), .ZN(new_n882));
  AOI211_X1 g0682(.A(KEYINPUT105), .B(new_n289), .C1(new_n882), .C2(new_n877), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n398), .B1(new_n885), .B2(new_n693), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n464), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n448), .A2(new_n453), .ZN(new_n889));
  INV_X1    g0689(.A(new_n693), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n448), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n398), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n465), .A2(new_n457), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n461), .A2(new_n462), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n464), .B1(new_n896), .B2(new_n386), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT81), .B1(new_n897), .B2(KEYINPUT18), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n399), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n289), .B1(new_n882), .B2(new_n877), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n385), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n896), .B1(new_n902), .B2(new_n883), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n890), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n894), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(new_n893), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n453), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n910), .A3(new_n398), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n904), .B1(new_n466), .B2(new_n399), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n426), .A2(new_n695), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n426), .A2(new_n918), .A3(new_n695), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n447), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n920), .B(new_n430), .C1(new_n446), .C2(new_n426), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n870), .B(new_n818), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT40), .B1(new_n915), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n889), .A2(new_n891), .A3(new_n398), .ZN(new_n927));
  INV_X1    g0727(.A(new_n892), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n929), .A2(new_n893), .ZN(new_n930));
  INV_X1    g0730(.A(new_n891), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n465), .A2(new_n651), .A3(new_n454), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n651), .B1(new_n465), .B2(new_n454), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n399), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n930), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n907), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n926), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n865), .B1(new_n872), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n872), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n934), .A2(new_n931), .ZN(new_n943));
  INV_X1    g0743(.A(new_n930), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n912), .A2(new_n913), .A3(new_n908), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n446), .A2(new_n426), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n695), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n907), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n653), .A2(new_n890), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n922), .A2(new_n923), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT102), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n695), .B(new_n816), .C1(new_n675), .C2(new_n684), .ZN(new_n955));
  INV_X1    g0755(.A(new_n813), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n827), .A2(KEYINPUT102), .A3(new_n813), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n952), .B1(new_n959), .B2(new_n915), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n667), .A2(new_n738), .A3(new_n750), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n666), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n864), .B1(new_n941), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n941), .ZN(new_n966));
  INV_X1    g0766(.A(new_n619), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(G116), .A3(new_n212), .A4(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT36), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n213), .A2(new_n308), .A3(new_n369), .A4(new_n370), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT101), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n972), .A2(new_n973), .B1(new_n296), .B2(G68), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n973), .B2(new_n972), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n688), .A3(new_n281), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n966), .A2(new_n971), .A3(new_n976), .ZN(G367));
  OR2_X1    g0777(.A1(new_n670), .A2(new_n671), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n978), .A2(new_n596), .A3(new_n706), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n596), .B(new_n672), .C1(new_n978), .C2(new_n706), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT108), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT43), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n743), .A2(new_n744), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n642), .A2(new_n706), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n989), .A2(new_n990), .B1(new_n740), .B2(new_n706), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n707), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT42), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(KEYINPUT42), .A3(new_n707), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n601), .B1(new_n992), .B2(new_n993), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n706), .B1(new_n1000), .B2(new_n633), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n988), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n994), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n705), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n999), .A2(new_n1001), .A3(new_n983), .A4(new_n985), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n713), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n708), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n994), .A2(KEYINPUT45), .A3(new_n708), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1004), .A2(KEYINPUT44), .A3(new_n1012), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n994), .B2(new_n708), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n705), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n704), .B1(new_n516), .B2(new_n706), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n707), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(new_n699), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n751), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1015), .A2(new_n1019), .A3(new_n705), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1021), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1010), .B1(new_n1029), .B2(new_n751), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1009), .B1(new_n1030), .B2(new_n754), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n779), .A2(new_n373), .B1(new_n772), .B2(new_n842), .ZN(new_n1032));
  INV_X1    g0832(.A(G143), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n793), .A2(new_n1033), .B1(new_n416), .B2(new_n777), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n760), .A2(new_n298), .B1(new_n768), .B2(new_n296), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G137), .B2(new_n765), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n246), .B1(new_n782), .B2(new_n308), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n772), .A2(new_n498), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT46), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n777), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G107), .A2(new_n1044), .B1(new_n771), .B2(G311), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n246), .B1(new_n848), .B2(G283), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n477), .A2(new_n478), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n761), .A2(new_n1048), .B1(new_n765), .B2(G317), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n782), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n778), .A2(G294), .B1(new_n1050), .B2(G97), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1046), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1041), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT47), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n758), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n232), .A2(new_n805), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n758), .B(new_n800), .C1(new_n712), .C2(new_n592), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n857), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1055), .B(new_n1058), .C1(new_n981), .C2(new_n809), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1031), .A2(new_n1059), .ZN(G387));
  OAI22_X1  g0860(.A1(new_n760), .A2(new_n296), .B1(new_n768), .B2(new_n416), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n251), .B(new_n1061), .C1(G150), .C2(new_n765), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n783), .A2(G97), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n778), .A2(new_n387), .B1(new_n773), .B2(G77), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n592), .A2(new_n1044), .B1(new_n771), .B2(G159), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n246), .B1(new_n765), .B2(G326), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n777), .A2(new_n832), .B1(new_n772), .B2(new_n775), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n761), .A2(G317), .B1(new_n848), .B2(new_n1048), .ZN(new_n1069));
  INV_X1    g0869(.A(G322), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n779), .B2(new_n767), .C1(new_n1070), .C2(new_n793), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1067), .B1(new_n498), .B2(new_n782), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n758), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n800), .B1(new_n702), .B2(new_n703), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n711), .A2(new_n802), .B1(new_n560), .B2(new_n712), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n711), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n300), .A2(G50), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT50), .ZN(new_n1088));
  AOI21_X1  g0888(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n264), .B2(new_n229), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT112), .B1(new_n1090), .B2(new_n805), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n857), .B1(new_n1094), .B2(new_n801), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1081), .A2(new_n1082), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT114), .B1(new_n1025), .B2(new_n751), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n713), .A3(new_n1026), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1025), .A2(new_n751), .A3(KEYINPUT114), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1096), .B1(new_n753), .B2(new_n1024), .C1(new_n1098), .C2(new_n1099), .ZN(G393));
  INV_X1    g0900(.A(new_n1028), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1026), .B1(new_n1101), .B2(new_n1020), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n1029), .A3(new_n713), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n793), .A2(new_n298), .B1(new_n373), .B2(new_n760), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n772), .A2(new_n416), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n777), .A2(new_n308), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G50), .C2(new_n778), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n246), .B1(new_n764), .B2(new_n1033), .C1(new_n300), .C2(new_n768), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AND4_X1   g0910(.A1(new_n837), .A2(new_n1105), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G317), .A2(new_n771), .B1(new_n761), .B2(G311), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n778), .A2(new_n1048), .B1(new_n773), .B2(G283), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n498), .B2(new_n777), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n251), .B1(new_n764), .B2(new_n1070), .C1(new_n775), .C2(new_n768), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1113), .A2(new_n786), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n758), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n240), .A2(new_n805), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n801), .C1(new_n494), .C2(new_n206), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n755), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1004), .B2(new_n800), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1101), .A2(new_n1020), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n754), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1103), .A2(new_n1124), .ZN(G390));
  XNOR2_X1  g0925(.A(new_n447), .B(new_n921), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n735), .B2(new_n818), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n870), .A2(G330), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n953), .A2(new_n1128), .A3(new_n816), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT102), .B1(new_n827), .B2(new_n813), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n695), .B1(new_n675), .B2(new_n684), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n954), .B(new_n956), .C1(new_n1131), .C2(new_n818), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1127), .A2(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n815), .A2(new_n654), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n695), .B(new_n1134), .C1(new_n745), .C2(new_n748), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT115), .B1(new_n1135), .B2(new_n956), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1134), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n749), .A2(new_n706), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT115), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n813), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT116), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n869), .ZN(new_n1143));
  OAI211_X1 g0943(.A(G330), .B(new_n818), .C1(new_n733), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1126), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1126), .A2(new_n735), .A3(new_n818), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n953), .A2(KEYINPUT116), .A3(new_n1144), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1141), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1133), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n467), .A2(new_n1128), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n962), .B(new_n1152), .C1(new_n661), .C2(new_n664), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1126), .B1(new_n1132), .B2(new_n1130), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n949), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n947), .A2(new_n950), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1136), .A2(new_n1126), .A3(new_n1140), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1159), .A2(new_n936), .A3(new_n1157), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1147), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1129), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n891), .B1(new_n653), .B2(new_n399), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n908), .B1(new_n1164), .B2(new_n930), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT39), .B1(new_n1165), .B2(new_n907), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n907), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n959), .B2(new_n949), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1159), .A2(new_n936), .A3(new_n1157), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1155), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1129), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1153), .B1(new_n1133), .B2(new_n1149), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1168), .A2(new_n1169), .A3(new_n1147), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n713), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n754), .A3(new_n1174), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n798), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n858), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n755), .B1(new_n387), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1044), .A2(G159), .B1(new_n848), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n850), .B2(new_n779), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT117), .Z(new_n1185));
  NOR2_X1   g0985(.A1(new_n772), .A2(new_n298), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT53), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n246), .B1(new_n760), .B2(new_n841), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G125), .B2(new_n765), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n771), .A2(G128), .B1(new_n1050), .B2(G50), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1107), .B1(G87), .B2(new_n773), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G107), .A2(new_n778), .B1(new_n771), .B2(G283), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n246), .B1(new_n765), .B2(G294), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n761), .A2(G116), .B1(new_n848), .B2(G97), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1185), .A2(new_n1191), .B1(new_n844), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1180), .B1(new_n1197), .B2(new_n758), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1178), .A2(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1177), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1176), .A2(new_n1200), .ZN(G378));
  NAND2_X1  g1001(.A1(new_n1175), .A2(new_n1154), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n915), .A2(new_n925), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n937), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n865), .B1(new_n936), .B2(new_n938), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n658), .A2(new_n660), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n305), .A2(new_n693), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1204), .A2(new_n1205), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n961), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n951), .A2(new_n960), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1214), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n936), .A2(new_n938), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(G330), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1221), .B2(new_n926), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1204), .A2(new_n1205), .A3(new_n1214), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1218), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1202), .A2(new_n1225), .A3(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n713), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1225), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n755), .B1(G50), .B2(new_n1179), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n251), .A2(new_n263), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n773), .B2(G77), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT118), .Z(new_n1233));
  AOI22_X1  g1033(.A1(new_n761), .A2(G107), .B1(new_n765), .B2(G283), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n311), .B2(new_n768), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n778), .A2(G97), .B1(new_n1050), .B2(G58), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n416), .B2(new_n777), .C1(new_n498), .C2(new_n793), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1233), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1231), .B(new_n296), .C1(G33), .C2(G41), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n773), .A2(new_n1182), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT119), .ZN(new_n1243));
  INV_X1    g1043(.A(G128), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n760), .A2(new_n1244), .B1(new_n768), .B2(new_n850), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G125), .B2(new_n771), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G150), .A2(new_n1044), .B1(new_n778), .B2(G132), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1050), .A2(G159), .ZN(new_n1251));
  AOI211_X1 g1051(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1241), .B1(KEYINPUT58), .B2(new_n1238), .C1(new_n1249), .C2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1230), .B1(new_n1254), .B2(new_n758), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1214), .B2(new_n799), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT120), .Z(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1225), .B2(new_n754), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1229), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(G375));
  INV_X1    g1061(.A(new_n1150), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1153), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1010), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1155), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n246), .B1(new_n783), .B2(G77), .ZN(new_n1266));
  XOR2_X1   g1066(.A(new_n1266), .B(KEYINPUT121), .Z(new_n1267));
  AOI22_X1  g1067(.A1(G107), .A2(new_n848), .B1(new_n765), .B2(G303), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n832), .B2(new_n760), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n779), .A2(new_n498), .B1(new_n311), .B2(new_n777), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n793), .A2(new_n775), .B1(new_n772), .B2(new_n494), .ZN(new_n1271));
  NOR4_X1   g1071(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n772), .A2(new_n373), .B1(new_n764), .B2(new_n1244), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT122), .Z(new_n1274));
  OAI221_X1 g1074(.A(new_n246), .B1(new_n768), .B2(new_n298), .C1(new_n850), .C2(new_n760), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n841), .A2(new_n793), .B1(new_n779), .B2(new_n1181), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n777), .A2(new_n296), .B1(new_n782), .B2(new_n842), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n758), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1279), .B(new_n755), .C1(G68), .C2(new_n1179), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n953), .B2(new_n798), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1150), .B2(new_n754), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1282), .ZN(G381));
  INV_X1    g1083(.A(KEYINPUT123), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G378), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1176), .A2(new_n1200), .A3(KEYINPUT123), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1260), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G390), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n862), .A3(new_n1289), .ZN(new_n1290));
  OR4_X1    g1090(.A1(G387), .A2(new_n1287), .A3(G381), .A4(new_n1290), .ZN(G407));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G343), .C2(new_n1287), .ZN(G409));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(new_n1289), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1031), .A2(new_n1059), .A3(G390), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G390), .B1(new_n1031), .B2(new_n1059), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1288), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1031), .A2(G390), .A3(new_n1059), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1295), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1217), .A2(new_n1224), .A3(KEYINPUT124), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT124), .B1(new_n1217), .B2(new_n1224), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n753), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1202), .A2(new_n1225), .A3(new_n1264), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1257), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1285), .B(new_n1286), .C1(new_n1307), .C2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G378), .B(new_n1258), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n694), .A2(G213), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1263), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1262), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n713), .A3(new_n1155), .A4(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(G384), .A3(new_n1282), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1318), .B2(new_n1282), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1313), .A2(new_n1314), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1303), .B1(new_n1304), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1314), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(G2897), .ZN(new_n1327));
  XOR2_X1   g1127(.A(new_n1327), .B(KEYINPUT125), .Z(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1321), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1328), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1319), .A3(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT126), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1323), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1335), .B1(new_n1336), .B2(KEYINPUT63), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1323), .A2(KEYINPUT126), .A3(new_n1304), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1324), .B(new_n1334), .C1(new_n1337), .C2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1326), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1340), .A2(KEYINPUT62), .A3(new_n1322), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT62), .B1(new_n1340), .B2(new_n1322), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1334), .B(KEYINPUT127), .C1(new_n1341), .C2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1303), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1323), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1340), .A2(KEYINPUT62), .A3(new_n1322), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT127), .B1(new_n1348), .B2(new_n1334), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1339), .B1(new_n1344), .B2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1312), .B1(new_n1260), .B2(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1322), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1303), .ZN(G402));
endmodule


