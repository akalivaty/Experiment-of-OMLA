//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  OAI21_X1  g0024(.A(KEYINPUT64), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n226), .A2(G1), .A3(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n209), .B1(new_n222), .B2(KEYINPUT1), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n218), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G50), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n225), .A2(new_n227), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n224), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n257), .A2(new_n225), .A3(new_n227), .A4(new_n254), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n223), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G68), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(G20), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(new_n266), .B(KEYINPUT12), .Z(new_n267));
  NAND3_X1  g0067(.A1(new_n230), .A2(G33), .A3(G77), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n268), .B1(new_n230), .B2(G68), .C1(new_n270), .C2(new_n202), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n225), .A2(new_n227), .A3(new_n254), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n267), .B1(KEYINPUT11), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n264), .B(new_n274), .C1(KEYINPUT11), .C2(new_n273), .ZN(new_n275));
  XOR2_X1   g0075(.A(new_n275), .B(KEYINPUT73), .Z(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n281), .A2(KEYINPUT69), .A3(G226), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n282), .B1(new_n279), .B2(new_n280), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G232), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n225), .A2(new_n227), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n223), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G238), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n296), .A2(new_n297), .B1(new_n298), .B2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT72), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g0103(.A(new_n299), .B(new_n302), .C1(new_n290), .C2(new_n291), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT71), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n301), .B2(KEYINPUT13), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n299), .B1(new_n290), .B2(new_n291), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n303), .B(new_n306), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n302), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G169), .B1(new_n316), .B2(new_n304), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT14), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(G169), .C1(new_n316), .C2(new_n304), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n276), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n316), .A2(new_n304), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n275), .B1(new_n324), .B2(G200), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n301), .A2(new_n307), .A3(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT71), .B1(new_n309), .B2(new_n310), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n328), .A2(G190), .A3(new_n303), .A4(new_n306), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G1698), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G222), .B1(G77), .B2(new_n335), .ZN(new_n337));
  INV_X1    g0137(.A(G223), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n281), .A2(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n291), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n295), .A2(new_n298), .ZN(new_n342));
  INV_X1    g0142(.A(new_n296), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(G226), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n345), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n224), .A2(new_n230), .A3(G1), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n272), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(G50), .A3(new_n263), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G50), .B2(new_n257), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n230), .A3(G33), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n255), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT9), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT10), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n345), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT67), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n341), .A2(new_n313), .A3(new_n344), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n230), .A3(G33), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n230), .B2(new_n372), .C1(new_n270), .C2(new_n353), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n272), .B1(new_n372), .B2(new_n349), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n262), .A2(G77), .A3(new_n263), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n336), .A2(G232), .B1(G107), .B2(new_n335), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n297), .B2(new_n339), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n291), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n342), .B1(new_n343), .B2(G244), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G179), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(G169), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n383), .A2(G200), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n382), .A2(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n377), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n332), .A2(new_n361), .A3(new_n368), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n281), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n265), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n217), .A2(new_n265), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n269), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT16), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n281), .A2(new_n393), .A3(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n335), .B2(new_n230), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(new_n400), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n272), .ZN(new_n409));
  OAI211_X1 g0209(.A(G223), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n410));
  OAI211_X1 g0210(.A(G226), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n278), .C2(new_n211), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n291), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n342), .B1(new_n343), .B2(G232), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n347), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(G200), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n354), .A2(new_n263), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n419), .A2(new_n259), .B1(new_n257), .B2(new_n354), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n409), .A2(new_n417), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT76), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n255), .B1(new_n401), .B2(new_n407), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n420), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(KEYINPUT76), .A3(new_n418), .A4(new_n417), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n409), .A2(new_n421), .A3(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n413), .A2(new_n414), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(G179), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n416), .A2(KEYINPUT74), .A3(new_n313), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n426), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT18), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT75), .B1(new_n435), .B2(new_n436), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT18), .B(new_n442), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n431), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n392), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n223), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n350), .A2(G87), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n369), .A2(new_n349), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT19), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n230), .B1(new_n287), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G87), .A2(G97), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n219), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n230), .B(G68), .C1(new_n333), .C2(new_n334), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n230), .A2(G33), .A3(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n453), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT80), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n272), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n454), .A2(new_n456), .B1(new_n453), .B2(new_n459), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT80), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n451), .B(new_n452), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G238), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n467));
  OAI211_X1 g0267(.A(G244), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n291), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n212), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n223), .A2(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n298), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n294), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G200), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n471), .A2(G190), .A3(new_n477), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n466), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT79), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n478), .B2(G179), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n350), .A2(new_n370), .A3(new_n450), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n452), .C1(new_n462), .C2(new_n464), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n471), .A2(KEYINPUT79), .A3(new_n313), .A4(new_n477), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n362), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n294), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT84), .B1(new_n494), .B2(new_n220), .ZN(new_n495));
  OAI211_X1 g0295(.A(G250), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n291), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n493), .A2(new_n501), .A3(G264), .A4(new_n294), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n495), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n492), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n475), .B1(new_n504), .B2(new_n490), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G274), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n347), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n495), .A2(new_n500), .A3(new_n506), .A4(new_n502), .ZN(new_n508));
  INV_X1    g0308(.A(G200), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n230), .A2(G107), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n256), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT25), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT83), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n350), .A2(G107), .A3(new_n450), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n281), .A2(new_n230), .A3(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n512), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n469), .A2(G20), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n230), .A2(KEYINPUT23), .A3(G107), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n523), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n281), .A2(new_n230), .A3(G87), .A4(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n524), .A2(new_n529), .A3(KEYINPUT24), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n272), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n531), .A3(new_n529), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n521), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n511), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n508), .A2(KEYINPUT85), .A3(G169), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n508), .A2(G169), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT85), .B1(new_n508), .B2(new_n313), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n489), .B(new_n539), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(new_n213), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n230), .B1(new_n372), .B2(new_n270), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n219), .B1(new_n394), .B2(new_n395), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n272), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n349), .A2(new_n213), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n350), .A2(G97), .A3(new_n450), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n506), .B1(new_n494), .B2(new_n214), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT4), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n557), .A2(KEYINPUT4), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G283), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n288), .B2(G250), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n313), .B(new_n555), .C1(new_n567), .C2(new_n291), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n563), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n556), .B2(new_n558), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n291), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n555), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n362), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n554), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT78), .B(new_n554), .C1(new_n568), .C2(new_n573), .ZN(new_n577));
  INV_X1    g0377(.A(new_n554), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n572), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n555), .B1(new_n567), .B2(new_n291), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n291), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n281), .A2(G257), .A3(new_n282), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n281), .A2(KEYINPUT81), .A3(G257), .A4(new_n282), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n288), .A2(G264), .B1(new_n335), .B2(G303), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G270), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n506), .B1(new_n494), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT21), .B(G169), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n594), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n339), .A2(new_n220), .B1(new_n597), .B2(new_n281), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  OAI211_X1 g0399(.A(G179), .B(new_n596), .C1(new_n599), .C2(new_n585), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n258), .A2(new_n261), .A3(G116), .A4(new_n450), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n278), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(G20), .B1(new_n604), .B2(new_n564), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n230), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n603), .B1(new_n608), .B2(new_n255), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n272), .B(KEYINPUT20), .C1(new_n605), .C2(new_n607), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n349), .A2(new_n606), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n602), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n601), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n509), .B1(new_n592), .B2(new_n594), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n347), .B(new_n596), .C1(new_n599), .C2(new_n585), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n596), .B1(new_n599), .B2(new_n585), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n613), .A3(G169), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n544), .A2(new_n584), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n449), .A2(new_n625), .ZN(G372));
  AND3_X1   g0426(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n542), .A2(new_n541), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n508), .A2(KEYINPUT85), .A3(G169), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n538), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n601), .A2(new_n613), .B1(new_n621), .B2(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n487), .B1(G179), .B2(new_n478), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n487), .B(KEYINPUT86), .C1(G179), .C2(new_n478), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n485), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(new_n480), .A3(new_n466), .A4(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n627), .A2(new_n633), .A3(new_n539), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n576), .A2(new_n577), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n489), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  INV_X1    g0447(.A(new_n574), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n642), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n643), .A2(new_n646), .A3(new_n638), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n449), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n368), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n435), .B(new_n436), .C1(new_n425), .C2(new_n420), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n323), .B1(new_n330), .B2(new_n386), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n424), .A2(new_n427), .B1(KEYINPUT17), .B2(new_n429), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n652), .B1(new_n658), .B2(new_n361), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n659), .ZN(G369));
  NAND2_X1  g0460(.A1(new_n256), .A2(new_n230), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  OAI21_X1  g0463(.A(G213), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G343), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n632), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n631), .B(new_n539), .C1(new_n538), .C2(new_n666), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n630), .A2(new_n667), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n631), .A2(new_n667), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT90), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n668), .B(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(new_n675), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n632), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n614), .A2(new_n623), .A3(new_n619), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n667), .A2(new_n613), .ZN(new_n686));
  MUX2_X1   g0486(.A(new_n684), .B(new_n685), .S(new_n686), .Z(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n673), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n683), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n207), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n455), .A2(new_n219), .A3(new_n606), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n234), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n644), .A2(new_n647), .A3(new_n489), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n638), .A2(new_n648), .A3(new_n641), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT26), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n643), .A2(new_n638), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n650), .A2(new_n666), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  INV_X1    g0507(.A(new_n478), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n581), .A2(new_n503), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT91), .B(new_n707), .C1(new_n709), .C2(new_n600), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n503), .A2(new_n708), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n592), .A2(new_n313), .A3(new_n594), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT30), .A4(new_n581), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n708), .A2(G179), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n620), .A3(new_n579), .A4(new_n508), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n710), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n711), .A2(new_n712), .A3(new_n581), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT91), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n666), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n519), .A2(new_n520), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n535), .A2(new_n536), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n533), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n510), .B2(new_n507), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n481), .A2(new_n488), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n630), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n627), .A2(new_n726), .A3(new_n685), .A4(new_n666), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n720), .B1(new_n727), .B2(KEYINPUT31), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n713), .A2(new_n715), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n717), .A2(new_n707), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n729), .B(new_n666), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(G330), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n706), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT92), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT92), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n699), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n224), .A2(G20), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n693), .A3(new_n223), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n687), .B2(G330), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n687), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n230), .A2(new_n347), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n313), .A2(new_n509), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  INV_X1    g0554(.A(G326), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n313), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G322), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n230), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n757), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n509), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(G303), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n230), .B1(new_n768), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G294), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n747), .A2(new_n760), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n281), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n764), .A2(new_n760), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(new_n768), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G283), .A2(new_n777), .B1(new_n779), .B2(G329), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n767), .A2(new_n771), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n769), .A2(new_n213), .ZN(new_n782));
  INV_X1    g0582(.A(new_n758), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n335), .B(new_n782), .C1(G58), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n766), .A2(G87), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n773), .A2(G68), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n777), .A2(G107), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n791), .B1(new_n372), .B2(new_n794), .C1(new_n202), .C2(new_n753), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n756), .A2(new_n781), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n229), .B1(G20), .B2(new_n362), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n745), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n281), .A2(new_n207), .ZN(new_n804));
  INV_X1    g0604(.A(G355), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(G116), .B2(new_n207), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n234), .A2(new_n472), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n249), .B2(new_n472), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n692), .A2(new_n281), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n801), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n798), .B1(new_n803), .B2(new_n810), .C1(new_n687), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n744), .A2(new_n812), .ZN(G396));
  OR2_X1    g0613(.A1(new_n797), .A2(new_n799), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n742), .B1(new_n814), .B2(G77), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  INV_X1    g0616(.A(new_n753), .ZN(new_n817));
  INV_X1    g0617(.A(new_n794), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n817), .A2(G303), .B1(new_n818), .B2(G116), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n281), .B(new_n782), .C1(G87), .C2(new_n777), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G283), .A2(new_n773), .B1(new_n783), .B2(G294), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G107), .A2(new_n766), .B1(new_n779), .B2(G311), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n776), .A2(new_n265), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G50), .B2(new_n766), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n281), .B1(new_n778), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G58), .B2(new_n770), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n758), .B1(new_n772), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n794), .A2(new_n789), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(G137), .C2(new_n817), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n826), .B(new_n829), .C1(new_n834), .C2(KEYINPUT34), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n823), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n816), .B1(new_n837), .B2(new_n797), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT101), .B1(new_n387), .B2(new_n666), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n376), .A2(new_n667), .A3(KEYINPUT100), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n377), .B2(new_n666), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n387), .A2(new_n390), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT101), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n386), .A2(new_n844), .A3(new_n667), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n839), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n838), .B1(new_n846), .B2(new_n800), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n705), .B(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n733), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n742), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n733), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n739), .A2(new_n223), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT107), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n665), .B1(new_n425), .B2(new_n420), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n448), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n429), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n653), .A2(new_n429), .A3(new_n859), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n858), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n861), .B2(new_n867), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n869), .B(new_n866), .C1(new_n448), .C2(new_n860), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT103), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n846), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n730), .A2(new_n710), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT31), .B(new_n667), .C1(new_n878), .C2(new_n718), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n729), .B1(new_n625), .B2(new_n666), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT106), .B(new_n879), .C1(new_n880), .C2(new_n720), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT106), .ZN(new_n882));
  INV_X1    g0682(.A(new_n879), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n728), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n877), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n320), .B(new_n318), .C1(new_n312), .C2(new_n313), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n276), .B(new_n667), .C1(new_n331), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n276), .A2(new_n667), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n322), .A2(new_n330), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT40), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n863), .A2(new_n864), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n865), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n860), .B1(new_n657), .B2(new_n654), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n894), .A2(new_n895), .B1(new_n864), .B2(new_n863), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n899), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n869), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n893), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n891), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n892), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n881), .A2(new_n884), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n449), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n857), .B(G330), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n876), .A2(new_n891), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n893), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G330), .A3(new_n907), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(G330), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n909), .A2(new_n911), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n322), .A2(new_n330), .A3(new_n888), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n888), .B1(new_n322), .B2(new_n330), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n650), .A2(new_n666), .A3(new_n846), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n386), .A2(new_n666), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n872), .B2(new_n875), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n654), .B1(new_n663), .B2(new_n664), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n905), .A2(new_n929), .A3(new_n871), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT39), .B1(new_n873), .B2(new_n874), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n322), .A2(new_n667), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n449), .B(new_n704), .C1(KEYINPUT29), .C2(new_n705), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n659), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n856), .B1(new_n919), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n919), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n234), .A2(new_n372), .A3(new_n397), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n265), .A2(G50), .ZN(new_n943));
  OAI211_X1 g0743(.A(G1), .B(new_n224), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n548), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n231), .B(G116), .C1(new_n945), .C2(KEYINPUT35), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(KEYINPUT35), .B2(new_n945), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT36), .Z(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n944), .A3(new_n948), .ZN(G367));
  OAI21_X1  g0749(.A(new_n627), .B1(new_n578), .B2(new_n666), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n648), .A2(new_n667), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n679), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT42), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(new_n631), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n666), .B1(new_n956), .B2(new_n644), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n666), .A2(new_n466), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n638), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n642), .B2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n955), .A2(new_n962), .A3(new_n961), .A4(new_n957), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n690), .A2(new_n953), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n693), .B(KEYINPUT41), .Z(new_n970));
  AOI21_X1  g0770(.A(new_n953), .B1(new_n676), .B2(new_n682), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n676), .A2(new_n682), .A3(new_n953), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n689), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n688), .B(new_n678), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n677), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n735), .B2(new_n736), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n974), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n682), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n952), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n972), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(new_n987), .A3(new_n690), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n976), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n970), .B1(new_n989), .B2(new_n737), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n741), .A2(new_n223), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n969), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n961), .A2(new_n801), .ZN(new_n994));
  INV_X1    g0794(.A(new_n809), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n244), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n996), .B(new_n803), .C1(new_n692), .C2(new_n370), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n745), .ZN(new_n998));
  INV_X1    g0798(.A(G294), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n335), .B1(new_n772), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G97), .A2(new_n777), .B1(new_n779), .B2(G317), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n597), .B2(new_n758), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G107), .C2(new_n770), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT46), .B1(new_n765), .B2(new_n606), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n606), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n818), .A2(G283), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n1006), .C1(new_n754), .C2(new_n762), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n770), .A2(G68), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n281), .C1(new_n217), .C2(new_n765), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n758), .A2(new_n831), .B1(new_n778), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n776), .A2(new_n372), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n772), .A2(new_n789), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n202), .B2(new_n794), .C1(new_n754), .C2(new_n830), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT47), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1007), .A2(KEYINPUT47), .A3(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n797), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n994), .B(new_n998), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n993), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT108), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT108), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n993), .A2(new_n1022), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(G387));
  NOR2_X1   g0825(.A1(new_n979), .A2(new_n694), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n978), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n737), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n673), .A2(new_n801), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n804), .A2(new_n696), .B1(G107), .B2(new_n207), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n240), .A2(G45), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n353), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G45), .B(new_n695), .C1(G68), .C2(G77), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n995), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1030), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n742), .B1(new_n1036), .B2(new_n803), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n202), .A2(new_n758), .B1(new_n772), .B2(new_n353), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n335), .B(new_n1038), .C1(G97), .C2(new_n777), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n817), .A2(G159), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n769), .A2(new_n369), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n761), .A2(new_n265), .B1(new_n778), .B2(new_n831), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n765), .A2(new_n372), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n281), .B1(new_n777), .B2(G116), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n773), .B1(new_n783), .B2(G317), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n597), .B2(new_n794), .C1(new_n754), .C2(new_n759), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n766), .A2(G294), .B1(new_n770), .B2(G283), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1047), .B1(new_n755), .B2(new_n778), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1046), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1037), .B1(new_n1058), .B2(new_n797), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1027), .A2(new_n992), .B1(new_n1029), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1028), .A2(new_n1060), .ZN(G393));
  INV_X1    g0861(.A(new_n979), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n988), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n690), .B1(new_n981), .B2(new_n987), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n693), .A3(new_n989), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n976), .A2(new_n988), .A3(new_n992), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n803), .B1(G97), .B2(new_n692), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n252), .A2(new_n809), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n745), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n797), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n817), .A2(G317), .B1(G311), .B2(new_n783), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n773), .B1(new_n779), .B2(G322), .ZN(new_n1074));
  INV_X1    g0874(.A(G283), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n765), .C1(new_n999), .C2(new_n761), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n787), .B(new_n335), .C1(new_n606), .C2(new_n769), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n753), .A2(new_n831), .B1(new_n789), .B2(new_n758), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n281), .B1(new_n769), .B2(new_n372), .C1(new_n211), .C2(new_n776), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G50), .A2(new_n773), .B1(new_n779), .B2(G143), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n265), .B2(new_n765), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(new_n354), .C2(new_n818), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1070), .B1(new_n1071), .B2(new_n1085), .C1(new_n952), .C2(new_n811), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1067), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1066), .A2(new_n1087), .ZN(G390));
  OAI211_X1 g0888(.A(new_n930), .B(new_n931), .C1(new_n925), .C2(new_n933), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n933), .B1(new_n905), .B2(new_n871), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n703), .A2(new_n666), .A3(new_n846), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1091), .A2(new_n924), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n890), .A2(KEYINPUT109), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT109), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n887), .A2(new_n889), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1090), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(G330), .B(new_n846), .C1(new_n728), .C2(new_n732), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(new_n922), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1089), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n910), .A2(G330), .A3(new_n846), .A4(new_n890), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT110), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT110), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n885), .A2(new_n1103), .A3(G330), .A4(new_n890), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1100), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n800), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n930), .A2(new_n931), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n742), .B1(new_n814), .B2(new_n354), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n785), .B(new_n335), .C1(new_n372), .C2(new_n769), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n758), .A2(new_n606), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n772), .A2(new_n219), .B1(new_n778), .B2(new_n999), .ZN(new_n1113));
  NOR4_X1   g0913(.A1(new_n1111), .A2(new_n824), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n213), .B2(new_n794), .C1(new_n1075), .C2(new_n753), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n753), .A2(new_n1116), .B1(new_n827), .B2(new_n758), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT115), .Z(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n772), .A2(new_n1010), .B1(new_n778), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n765), .A2(new_n831), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1121), .A2(new_n1122), .B1(new_n789), .B2(new_n769), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1120), .B(new_n1123), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n281), .B1(new_n776), .B2(new_n202), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT113), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n818), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1124), .A2(new_n1126), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1115), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1110), .B1(new_n1132), .B2(new_n797), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1107), .A2(new_n992), .B1(new_n1109), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1100), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1092), .B1(new_n922), .B2(new_n1098), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n885), .A2(G330), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n1096), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1098), .A2(new_n922), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1102), .A2(new_n1104), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n923), .A2(new_n924), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n938), .A2(new_n916), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1137), .A2(new_n1144), .A3(KEYINPUT111), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT111), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1140), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1147), .B1(new_n1150), .B2(new_n1107), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT112), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1150), .B2(new_n1107), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1137), .B(KEYINPUT112), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n693), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1134), .B1(new_n1152), .B2(new_n1156), .ZN(G378));
  NAND2_X1  g0957(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1145), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1107), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT111), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1150), .A2(new_n1147), .A3(new_n1107), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n361), .A2(new_n368), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n665), .B1(new_n352), .B2(new_n357), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n928), .B2(new_n935), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n934), .A3(new_n927), .A4(new_n926), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(G330), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n892), .A2(new_n908), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n915), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1163), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1159), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1177), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n694), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1168), .A2(new_n1108), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n742), .B1(new_n814), .B2(G50), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n281), .A2(G41), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n779), .A2(G283), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n217), .B2(new_n776), .C1(new_n369), .C2(new_n761), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1187), .A2(new_n1044), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G97), .A2(new_n773), .B1(new_n783), .B2(G107), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1008), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(G116), .C2(new_n817), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1188), .B1(new_n1194), .B2(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(KEYINPUT58), .B2(new_n1194), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n777), .C2(G159), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT118), .B(G124), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n753), .A2(new_n1119), .B1(new_n831), .B2(new_n769), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT117), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n783), .A2(G128), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n761), .B2(new_n1010), .C1(new_n827), .C2(new_n772), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n766), .B2(new_n1128), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1197), .B1(new_n778), .B2(new_n1198), .C1(new_n1204), .C2(KEYINPUT59), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1196), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1185), .B1(new_n1207), .B2(new_n797), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1177), .A2(new_n992), .B1(new_n1184), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT119), .B1(new_n1183), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1183), .A2(KEYINPUT119), .A3(new_n1210), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1158), .A2(new_n992), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1096), .A2(new_n799), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G97), .A2(new_n766), .B1(new_n779), .B2(G303), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n606), .B2(new_n772), .C1(new_n1075), .C2(new_n758), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1218), .A2(new_n281), .A3(new_n1012), .A4(new_n1041), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n817), .A2(G294), .B1(new_n818), .B2(G107), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n281), .B1(new_n769), .B2(new_n202), .C1(new_n217), .C2(new_n776), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n761), .A2(new_n831), .B1(new_n778), .B2(new_n1116), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1010), .A2(new_n758), .B1(new_n765), .B2(new_n789), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n817), .A2(G132), .B1(new_n773), .B2(new_n1128), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1219), .A2(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n742), .B1(G68), .B2(new_n814), .C1(new_n1226), .C2(new_n1071), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT120), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1216), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1215), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1150), .A2(new_n970), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1230), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G381));
  NAND2_X1  g1035(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1210), .B1(new_n1236), .B2(new_n693), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT119), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G378), .B1(new_n1239), .B2(new_n1211), .ZN(new_n1240));
  OR2_X1    g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1241), .A2(G384), .A3(G390), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n1024), .A3(new_n1234), .A4(new_n1242), .ZN(G407));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1021), .A2(new_n1023), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1241), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n993), .A2(G390), .A3(new_n1019), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n993), .A2(G390), .A3(new_n1253), .A4(new_n1019), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1248), .A2(new_n1250), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(KEYINPUT123), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n993), .A2(G390), .A3(new_n1257), .A4(new_n1019), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1020), .A2(new_n1247), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1250), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1255), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  OAI21_X1  g1066(.A(G378), .B1(new_n1183), .B2(new_n1210), .ZN(new_n1267));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1209), .B(new_n1134), .C1(new_n1152), .C2(new_n1156), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1163), .A2(new_n970), .A3(new_n1178), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT121), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1144), .A2(KEYINPUT121), .A3(KEYINPUT60), .A4(new_n1145), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n693), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT60), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1230), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1230), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1283), .B1(new_n1286), .B2(KEYINPUT122), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT122), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1282), .A2(new_n1288), .A3(G384), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1267), .A2(new_n1273), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1267), .A2(new_n1273), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1266), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1267), .A2(new_n1273), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1269), .A2(G2897), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1286), .A2(KEYINPUT122), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1288), .B1(new_n1282), .B2(G384), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1299), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1283), .A4(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1297), .B1(new_n1298), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1264), .B1(new_n1296), .B2(new_n1306), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1267), .A2(new_n1273), .B1(new_n1300), .B2(new_n1304), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1291), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1273), .A4(new_n1290), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1311), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1307), .B1(new_n1315), .B2(new_n1316), .ZN(G405));
  NAND3_X1  g1117(.A1(new_n1245), .A2(new_n1267), .A3(new_n1263), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1267), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1264), .B1(new_n1240), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1290), .A2(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1318), .A2(new_n1320), .A3(KEYINPUT127), .A4(new_n1290), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(G402));
endmodule


