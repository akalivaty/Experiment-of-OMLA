//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT66), .A2(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G119), .A3(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT67), .B1(new_n191), .B2(G119), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n199), .A3(G119), .A4(new_n193), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n197), .B2(new_n200), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n198), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT66), .A2(G116), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT66), .A2(G116), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n195), .B1(new_n207), .B2(G119), .ZN(new_n208));
  INV_X1    g022(.A(new_n200), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT64), .A3(G143), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n218), .B2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(G128), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(G137), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n231), .A2(G137), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n233), .A2(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n225), .A2(new_n244), .B1(new_n245), .B2(new_n242), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n237), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n229), .A2(new_n241), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT28), .B1(new_n213), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n201), .A2(new_n202), .A3(new_n189), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n210), .B2(new_n211), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n237), .A2(new_n240), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT69), .B1(new_n228), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n214), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n217), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(new_n221), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n241), .B(new_n259), .C1(new_n263), .C2(new_n220), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n249), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n253), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n213), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n228), .B2(new_n257), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n241), .B(new_n271), .C1(new_n263), .C2(new_n220), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n272), .A3(new_n265), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n267), .A2(new_n269), .B1(new_n256), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n252), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n277), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G101), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n267), .A2(new_n269), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n273), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n258), .A2(new_n264), .A3(KEYINPUT30), .A4(new_n265), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n256), .A3(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n284), .A2(new_n288), .A3(new_n282), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n276), .A2(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n256), .A2(new_n266), .A3(new_n253), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT70), .B1(new_n268), .B2(new_n213), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n288), .B(new_n282), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n284), .A2(KEYINPUT72), .A3(new_n288), .A4(new_n282), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(KEYINPUT31), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n188), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n282), .B(new_n252), .C1(new_n274), .C2(new_n275), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n301), .B2(new_n283), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n267), .A2(new_n269), .B1(new_n256), .B2(new_n266), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n252), .B(new_n304), .C1(new_n305), .C2(new_n275), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n256), .A2(new_n266), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n292), .B2(new_n293), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n252), .A4(new_n304), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n303), .A2(new_n307), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n299), .A2(KEYINPUT32), .B1(new_n314), .B2(G472), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n299), .B2(KEYINPUT32), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n276), .A2(new_n283), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n284), .A2(new_n290), .A3(new_n288), .A4(new_n282), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n298), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n187), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT32), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT73), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G475), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT77), .A2(G125), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(G125), .A2(G140), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT90), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(KEYINPUT77), .A2(G125), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT77), .A2(G125), .ZN(new_n335));
  OAI21_X1  g149(.A(G140), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n337));
  INV_X1    g151(.A(new_n332), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G146), .ZN(new_n342));
  INV_X1    g156(.A(G237), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G214), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n218), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT18), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n235), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n346), .A2(KEYINPUT18), .A3(G131), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n216), .B1(new_n333), .B2(new_n339), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n216), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT91), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n342), .B(new_n352), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n329), .A2(new_n330), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n332), .B1(new_n358), .B2(G140), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT16), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n326), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n216), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI221_X1 g179(.A(G146), .B1(new_n362), .B2(new_n363), .C1(new_n359), .C2(new_n360), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n348), .A2(KEYINPUT17), .A3(G131), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n348), .A2(G131), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT17), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n346), .A2(new_n235), .A3(new_n347), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n365), .A2(new_n366), .A3(new_n367), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n374), .B(G104), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n357), .A2(new_n372), .A3(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n325), .B1(new_n379), .B2(new_n313), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT19), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT92), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n354), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(KEYINPUT19), .C1(new_n382), .C2(new_n383), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(new_n216), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n361), .A2(new_n216), .A3(new_n364), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n368), .A2(new_n370), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n353), .A2(new_n356), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n353), .A2(new_n341), .B1(new_n351), .B2(new_n350), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n390), .A2(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n378), .B1(new_n396), .B2(new_n375), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n397), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n381), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G952), .ZN(new_n403));
  AOI211_X1 g217(.A(G953), .B(new_n403), .C1(G234), .C2(G237), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT21), .B(G898), .Z(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT96), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n313), .B(new_n344), .C1(G234), .C2(G237), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(G217), .A3(new_n344), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n218), .A2(G128), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n214), .A2(G143), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n231), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n419), .A3(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n417), .B1(new_n214), .B2(G143), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT93), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n416), .B1(new_n423), .B2(new_n231), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n192), .A2(G122), .A3(new_n193), .ZN(new_n425));
  INV_X1    g239(.A(G107), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n191), .A2(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n425), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT94), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G107), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n218), .A2(G128), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n214), .A2(G143), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(KEYINPUT13), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n421), .A2(KEYINPUT93), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n419), .B1(new_n414), .B2(new_n417), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G134), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n436), .A2(new_n443), .A3(new_n444), .A4(new_n416), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n432), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .A4(new_n193), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n427), .B1(new_n207), .B2(G122), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n416), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n231), .B1(new_n414), .B2(new_n415), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n435), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n413), .B1(new_n446), .B2(new_n456), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n412), .B(new_n455), .C1(new_n432), .C2(new_n445), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT95), .B(new_n313), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G478), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT15), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n424), .A2(new_n431), .A3(KEYINPUT94), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n452), .B1(new_n442), .B2(G134), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n444), .B1(new_n464), .B2(new_n436), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n456), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n412), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n455), .B1(new_n432), .B2(new_n445), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n413), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n461), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(KEYINPUT95), .A3(new_n313), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n402), .A2(new_n409), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G221), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n411), .B2(new_n313), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n344), .A2(G227), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n478), .B(new_n479), .Z(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n228), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(KEYINPUT82), .A2(G104), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n426), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT82), .A2(G104), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G101), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n426), .A3(G104), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT3), .A2(G107), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n483), .A2(new_n426), .A3(new_n486), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(G104), .B2(G107), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n260), .B2(new_n245), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n482), .A2(new_n496), .B1(new_n499), .B2(new_n481), .ZN(new_n500));
  INV_X1    g314(.A(new_n249), .ZN(new_n501));
  INV_X1    g315(.A(new_n487), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n489), .A2(new_n490), .ZN(new_n503));
  OAI21_X1  g317(.A(G101), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(G101), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n246), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n500), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n501), .B1(new_n500), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n480), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n495), .A2(new_n228), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n499), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n249), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT12), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n500), .A2(new_n501), .A3(new_n508), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n520), .A3(new_n516), .ZN(new_n521));
  INV_X1    g335(.A(new_n480), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT85), .B(G469), .Z(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT12), .B(new_n515), .C1(new_n499), .C2(new_n512), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n520), .B1(new_n513), .B2(new_n516), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n509), .A2(new_n510), .A3(new_n480), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT84), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n480), .ZN(new_n534));
  INV_X1    g348(.A(new_n510), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n519), .A3(new_n522), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G469), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n526), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n474), .A2(new_n477), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT5), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n197), .B2(new_n200), .ZN(new_n546));
  INV_X1    g360(.A(G119), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n547), .A3(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G113), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n544), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT5), .B1(new_n208), .B2(new_n209), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT86), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n495), .A2(new_n202), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT87), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n203), .A2(new_n212), .A3(new_n507), .A4(new_n505), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT87), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G122), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n556), .A2(new_n561), .A3(new_n557), .A4(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n566), .A3(new_n562), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n246), .A2(new_n362), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n228), .A2(KEYINPUT88), .A3(new_n362), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT88), .B1(new_n228), .B2(new_n362), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G224), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G953), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n565), .A2(new_n567), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n554), .B1(new_n546), .B2(new_n549), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n550), .A2(new_n553), .A3(new_n210), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(new_n496), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n561), .B(KEYINPUT8), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT89), .B1(new_n570), .B2(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n228), .A2(new_n362), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n569), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n587), .A3(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT7), .B1(new_n573), .B2(G953), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n572), .A2(new_n589), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n590), .A3(new_n564), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n313), .ZN(new_n593));
  OAI21_X1  g407(.A(G210), .B1(G237), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n576), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n593), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n565), .A2(new_n567), .A3(new_n575), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n543), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n542), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G217), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(G234), .B2(new_n313), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n365), .A2(new_n366), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n547), .A2(G128), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n547), .A2(G128), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(KEYINPUT23), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G110), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n611), .A2(KEYINPUT76), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT24), .B(G110), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(KEYINPUT75), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(KEYINPUT75), .ZN(new_n615));
  INV_X1    g429(.A(new_n609), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n608), .ZN(new_n617));
  OR3_X1    g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(KEYINPUT76), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n606), .A2(new_n612), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n610), .A2(G110), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n621), .A2(new_n622), .B1(new_n216), .B2(new_n354), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n623), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT78), .B1(new_n623), .B2(new_n366), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT22), .B(G137), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n344), .A2(G221), .A3(G234), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n366), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT78), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n623), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n620), .A3(new_n629), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT80), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT80), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n603), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT79), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT25), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n631), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n648), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n631), .A2(new_n637), .A3(new_n650), .A4(new_n646), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n605), .A2(new_n642), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n324), .A2(new_n601), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G101), .ZN(G3));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n468), .B2(new_n413), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(KEYINPUT33), .C1(new_n458), .C2(new_n457), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n467), .B(new_n469), .C1(new_n655), .C2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n659), .A3(G478), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n460), .A2(new_n313), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n467), .B2(new_n469), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n460), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n402), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n543), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n595), .B1(new_n576), .B2(new_n593), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n597), .A2(new_n598), .A3(new_n594), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n409), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(G902), .B1(new_n291), .B2(new_n298), .ZN(new_n676));
  INV_X1    g490(.A(G472), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n321), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n652), .A2(new_n541), .A3(new_n477), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT99), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT34), .B(G104), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  AND3_X1   g498(.A1(new_n357), .A2(new_n375), .A3(new_n372), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n389), .A2(new_n387), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n388), .B1(new_n340), .B2(KEYINPUT19), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(G146), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n391), .A2(new_n392), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n357), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n685), .B1(new_n690), .B2(new_n376), .ZN(new_n691));
  INV_X1    g505(.A(new_n399), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT20), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n380), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n473), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n674), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n680), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT35), .B(G107), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G9));
  NOR2_X1   g514(.A1(new_n630), .A2(KEYINPUT36), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n626), .B(new_n701), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n649), .A2(new_n651), .B1(new_n605), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n678), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n601), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  NAND2_X1  g521(.A1(new_n647), .A2(new_n648), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n603), .A3(new_n651), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n702), .A2(new_n605), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n541), .A2(new_n477), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n408), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n404), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n695), .A2(new_n473), .A3(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n600), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n324), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  NAND2_X1  g534(.A1(new_n309), .A2(new_n283), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n296), .A2(new_n297), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n677), .B1(new_n722), .B2(new_n313), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n299), .B2(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n317), .A2(new_n323), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(KEYINPUT100), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(KEYINPUT100), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n596), .A2(new_n599), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT38), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT38), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n716), .B(KEYINPUT39), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n541), .A2(new_n477), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n737));
  INV_X1    g551(.A(new_n473), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n695), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n543), .A3(new_n703), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n736), .B2(KEYINPUT40), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n729), .A2(new_n734), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT101), .B(G143), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G45));
  INV_X1    g558(.A(new_n716), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n695), .A2(new_n664), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n477), .A3(new_n541), .A4(new_n711), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n600), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n324), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT102), .B(G146), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G48));
  AND2_X1   g565(.A1(new_n524), .A2(new_n525), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n524), .A2(new_n540), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n476), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n675), .A2(new_n324), .A3(new_n652), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND4_X1  g573(.A1(new_n697), .A2(new_n324), .A3(new_n652), .A4(new_n756), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AND2_X1   g575(.A1(new_n756), .A2(new_n672), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n324), .A2(new_n762), .A3(new_n474), .A4(new_n711), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  AOI21_X1  g578(.A(new_n677), .B1(new_n320), .B2(new_n313), .ZN(new_n765));
  INV_X1    g579(.A(new_n652), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n252), .B1(new_n305), .B2(new_n275), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n767), .A2(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n188), .B1(new_n768), .B2(new_n298), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n739), .B(new_n543), .C1(new_n596), .C2(new_n599), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n772), .A3(new_n673), .A4(new_n756), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT103), .B(G122), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G24));
  NAND3_X1  g589(.A1(new_n665), .A2(new_n402), .A3(new_n716), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n765), .A2(new_n776), .A3(new_n769), .A4(new_n703), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n762), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  NAND2_X1  g593(.A1(new_n321), .A2(new_n322), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n314), .A2(G472), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n540), .A2(new_n313), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n524), .B2(new_n525), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n534), .A2(KEYINPUT104), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n533), .A2(new_n787), .A3(new_n480), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(G469), .A3(new_n536), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n476), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n670), .A2(new_n790), .A3(new_n543), .A4(new_n671), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n776), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(new_n792), .A3(new_n652), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT42), .ZN(new_n794));
  INV_X1    g608(.A(new_n791), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n324), .A2(new_n652), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n235), .ZN(G33));
  INV_X1    g613(.A(new_n717), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n324), .A2(new_n652), .A3(new_n800), .A4(new_n795), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND4_X1  g616(.A1(new_n786), .A2(KEYINPUT45), .A3(new_n536), .A4(new_n788), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n532), .A2(new_n538), .ZN(new_n804));
  OAI211_X1 g618(.A(G469), .B(new_n803), .C1(new_n804), .C2(KEYINPUT45), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT105), .Z(new_n806));
  INV_X1    g620(.A(new_n784), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT46), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(KEYINPUT106), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n808), .B2(KEYINPUT46), .ZN(new_n812));
  OAI221_X1 g626(.A(new_n526), .B1(KEYINPUT46), .B2(new_n808), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n477), .A3(new_n735), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n670), .A2(new_n543), .A3(new_n671), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n402), .A2(new_n664), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT43), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n678), .A3(new_n711), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n814), .B(new_n820), .C1(new_n819), .C2(new_n818), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  NOR2_X1   g636(.A1(new_n810), .A2(new_n812), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n526), .B1(new_n808), .B2(KEYINPUT46), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT107), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n825), .A2(new_n476), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n813), .B(new_n477), .C1(new_n827), .C2(new_n828), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n324), .A2(new_n652), .A3(new_n776), .A4(new_n815), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  NAND3_X1  g648(.A1(new_n652), .A2(new_n543), .A3(new_n477), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n816), .B1(new_n835), .B2(KEYINPUT108), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(KEYINPUT108), .B2(new_n835), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT109), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n754), .B(KEYINPUT49), .Z(new_n839));
  OR4_X1    g653(.A1(new_n729), .A2(new_n838), .A3(new_n734), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n770), .A2(new_n404), .A3(new_n817), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n756), .A2(new_n672), .ZN(new_n842));
  OAI211_X1 g656(.A(G952), .B(new_n344), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n817), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n756), .A2(new_n730), .A3(new_n543), .A4(new_n404), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n652), .A3(new_n783), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT48), .Z(new_n848));
  INV_X1    g662(.A(new_n668), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n729), .A2(new_n766), .A3(new_n845), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n843), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(new_n695), .A3(new_n664), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n733), .A2(new_n669), .A3(new_n756), .ZN(new_n853));
  OR4_X1    g667(.A1(KEYINPUT117), .A2(new_n853), .A3(KEYINPUT50), .A4(new_n841), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n853), .B2(new_n841), .ZN(new_n856));
  INV_X1    g670(.A(new_n298), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n251), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n319), .B1(new_n858), .B2(new_n282), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n187), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n711), .C1(new_n676), .C2(new_n677), .ZN(new_n861));
  INV_X1    g675(.A(new_n846), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n854), .B(new_n856), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n755), .A2(new_n477), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n830), .B2(new_n831), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n841), .A2(new_n815), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n851), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT110), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n462), .A2(new_n472), .A3(new_n716), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n402), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n462), .A2(new_n472), .A3(new_n716), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT110), .B1(new_n695), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n712), .A3(new_n815), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT111), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(new_n324), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n878), .B2(new_n324), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT112), .B1(new_n777), .B2(new_n795), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n861), .A2(new_n791), .A3(new_n884), .A4(new_n776), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n801), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n882), .A2(new_n886), .A3(new_n798), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n703), .A2(new_n790), .A3(new_n716), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n771), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n725), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n719), .A2(new_n749), .A3(new_n778), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n324), .B1(new_n718), .B2(new_n748), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(KEYINPUT52), .A3(new_n778), .A4(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n666), .A2(new_n696), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n672), .A2(new_n673), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n680), .A2(new_n898), .B1(new_n601), .B2(new_n704), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n653), .A3(new_n763), .A4(new_n773), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n757), .A2(new_n760), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n887), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n891), .A2(KEYINPUT113), .A3(new_n892), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT113), .B(KEYINPUT114), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n895), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n895), .ZN(new_n908));
  INV_X1    g722(.A(new_n906), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n904), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  MUX2_X1   g726(.A(new_n903), .B(new_n911), .S(new_n912), .Z(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n913), .A2(KEYINPUT115), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT115), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n907), .A4(new_n910), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n903), .A2(new_n918), .A3(new_n912), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n903), .B2(new_n912), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n914), .B(new_n917), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n869), .A2(new_n923), .A3(new_n870), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n869), .A2(new_n870), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT118), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n871), .B(new_n922), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n840), .B1(new_n927), .B2(new_n928), .ZN(G75));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n565), .A2(new_n567), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n575), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  AND2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n934), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n344), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  NAND2_X1  g755(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n921), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n931), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n784), .B(KEYINPUT57), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT120), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n944), .A2(new_n949), .A3(new_n945), .A4(new_n946), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n511), .A2(new_n523), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT121), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n932), .A2(new_n806), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n948), .B2(new_n950), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n940), .B1(new_n954), .B2(new_n958), .ZN(G54));
  NAND4_X1  g773(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n691), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n691), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n940), .ZN(G60));
  NAND2_X1  g777(.A1(new_n657), .A2(new_n659), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n661), .B(KEYINPUT59), .Z(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n922), .B2(new_n965), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n964), .A2(new_n944), .A3(new_n945), .A4(new_n965), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n940), .A3(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT122), .Z(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n931), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n642), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n940), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n702), .B(KEYINPUT123), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT61), .Z(G66));
  NOR2_X1   g791(.A1(new_n902), .A2(G953), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT124), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n407), .B2(new_n573), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n935), .B1(G898), .B2(new_n344), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT126), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n981), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n286), .A2(new_n287), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n686), .A2(new_n687), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(new_n988));
  NAND2_X1  g802(.A1(G900), .A2(G953), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n814), .A2(new_n652), .A3(new_n772), .A4(new_n783), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n894), .A2(new_n778), .A3(new_n801), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(new_n798), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n821), .A2(new_n990), .A3(new_n833), .A4(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n988), .B(new_n989), .C1(new_n993), .C2(G953), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n742), .A2(new_n778), .A3(new_n894), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT62), .Z(new_n996));
  AOI211_X1 g810(.A(new_n815), .B(new_n736), .C1(new_n666), .C2(new_n696), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n324), .A3(new_n652), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n821), .A2(new_n833), .A3(new_n996), .A4(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n999), .A2(new_n344), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n994), .B1(new_n1000), .B2(new_n988), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n344), .B1(G227), .B2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(new_n301), .A2(new_n282), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  INV_X1    g820(.A(new_n902), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1008), .A2(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(KEYINPUT127), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1004), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1006), .B1(new_n993), .B2(new_n1007), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n301), .A2(new_n282), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n940), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n296), .A2(new_n297), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n282), .B1(new_n284), .B2(new_n288), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1006), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1014), .B1(new_n913), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1011), .A2(new_n1018), .ZN(G57));
endmodule


