

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765;

  BUF_X1 U374 ( .A(n725), .Z(n729) );
  INV_X1 U375 ( .A(G128), .ZN(n438) );
  NOR2_X2 U376 ( .A1(G953), .A2(G237), .ZN(n446) );
  INV_X4 U377 ( .A(G953), .ZN(n744) );
  NOR2_X1 U378 ( .A1(n641), .A2(n733), .ZN(n643) );
  NOR2_X1 U379 ( .A1(n653), .A2(n733), .ZN(n654) );
  AND2_X1 U380 ( .A1(n696), .A2(n521), .ZN(n605) );
  XNOR2_X2 U381 ( .A(G113), .B(KEYINPUT3), .ZN(n387) );
  XNOR2_X2 U382 ( .A(n487), .B(G134), .ZN(n443) );
  BUF_X1 U383 ( .A(n631), .Z(n734) );
  NAND2_X1 U384 ( .A1(n383), .A2(n583), .ZN(n753) );
  NAND2_X1 U385 ( .A1(n600), .A2(n547), .ZN(n393) );
  OR2_X1 U386 ( .A1(n684), .A2(n683), .ZN(n689) );
  BUF_X1 U387 ( .A(n521), .Z(n695) );
  BUF_X1 U388 ( .A(n518), .Z(n407) );
  XNOR2_X1 U389 ( .A(n479), .B(KEYINPUT10), .ZN(n750) );
  AND2_X2 U390 ( .A1(n636), .A2(n635), .ZN(n725) );
  XNOR2_X2 U391 ( .A(n439), .B(n438), .ZN(n487) );
  XNOR2_X2 U392 ( .A(n474), .B(n473), .ZN(n741) );
  XNOR2_X2 U393 ( .A(n445), .B(n444), .ZN(n474) );
  AND2_X1 U394 ( .A1(n578), .A2(n579), .ZN(n385) );
  XNOR2_X1 U395 ( .A(n387), .B(G119), .ZN(n445) );
  AND2_X1 U396 ( .A1(n577), .A2(n763), .ZN(n578) );
  XNOR2_X1 U397 ( .A(n443), .B(n442), .ZN(n461) );
  XNOR2_X1 U398 ( .A(n609), .B(KEYINPUT1), .ZN(n521) );
  XNOR2_X1 U399 ( .A(n384), .B(n580), .ZN(n383) );
  XNOR2_X1 U400 ( .A(n398), .B(n380), .ZN(n379) );
  XNOR2_X1 U401 ( .A(n381), .B(n353), .ZN(n380) );
  NAND2_X1 U402 ( .A1(n364), .A2(n375), .ZN(n373) );
  INV_X1 U403 ( .A(n559), .ZN(n364) );
  INV_X1 U404 ( .A(KEYINPUT40), .ZN(n367) );
  NAND2_X1 U405 ( .A1(n370), .A2(KEYINPUT40), .ZN(n369) );
  NAND2_X1 U406 ( .A1(n373), .A2(n372), .ZN(n370) );
  INV_X1 U407 ( .A(n376), .ZN(n374) );
  NAND2_X1 U408 ( .A1(n725), .A2(G210), .ZN(n392) );
  AND2_X1 U409 ( .A1(n595), .A2(n584), .ZN(n591) );
  XNOR2_X1 U410 ( .A(n396), .B(n382), .ZN(n381) );
  INV_X1 U411 ( .A(KEYINPUT85), .ZN(n382) );
  XNOR2_X1 U412 ( .A(G137), .B(G128), .ZN(n396) );
  XNOR2_X1 U413 ( .A(n524), .B(n523), .ZN(n682) );
  OR2_X1 U414 ( .A1(n637), .A2(G902), .ZN(n454) );
  AND2_X1 U415 ( .A1(n686), .A2(n500), .ZN(n501) );
  OR2_X1 U416 ( .A1(n518), .A2(n698), .ZN(n520) );
  OR2_X1 U417 ( .A1(n650), .A2(G902), .ZN(n469) );
  XNOR2_X1 U418 ( .A(n461), .B(n394), .ZN(n752) );
  XNOR2_X1 U419 ( .A(n741), .B(n475), .ZN(n493) );
  BUF_X1 U420 ( .A(n682), .Z(n715) );
  XNOR2_X1 U421 ( .A(n399), .B(n379), .ZN(n400) );
  NAND2_X1 U422 ( .A1(n725), .A2(G475), .ZN(n363) );
  NAND2_X1 U423 ( .A1(n374), .A2(n373), .ZN(n545) );
  NAND2_X1 U424 ( .A1(n368), .A2(n365), .ZN(n557) );
  NAND2_X1 U425 ( .A1(n374), .A2(n355), .ZN(n365) );
  AND2_X1 U426 ( .A1(n371), .A2(n369), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n576), .B(KEYINPUT112), .ZN(n763) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(G60) );
  INV_X1 U429 ( .A(KEYINPUT60), .ZN(n359) );
  NAND2_X1 U430 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n363), .B(n358), .ZN(n362) );
  INV_X1 U432 ( .A(KEYINPUT56), .ZN(n388) );
  XNOR2_X1 U433 ( .A(n392), .B(n391), .ZN(n390) );
  XOR2_X1 U434 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n353) );
  XOR2_X1 U435 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n354) );
  AND2_X1 U436 ( .A1(n373), .A2(n366), .ZN(n355) );
  AND2_X1 U437 ( .A1(n609), .A2(n538), .ZN(n356) );
  XOR2_X1 U438 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n357) );
  INV_X1 U439 ( .A(n669), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n493), .B(n492), .ZN(n721) );
  XNOR2_X1 U441 ( .A(n728), .B(n727), .ZN(n358) );
  INV_X1 U442 ( .A(n733), .ZN(n361) );
  AND2_X1 U443 ( .A1(n372), .A2(n367), .ZN(n366) );
  NAND2_X1 U444 ( .A1(n376), .A2(KEYINPUT40), .ZN(n371) );
  NOR2_X1 U445 ( .A1(n684), .A2(n357), .ZN(n375) );
  NAND2_X1 U446 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U447 ( .A1(n684), .A2(n357), .ZN(n377) );
  NAND2_X1 U448 ( .A1(n559), .A2(n357), .ZN(n378) );
  NAND2_X1 U449 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n558), .B(KEYINPUT46), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(G51) );
  NAND2_X1 U452 ( .A1(n390), .A2(n361), .ZN(n389) );
  INV_X1 U453 ( .A(n724), .ZN(n391) );
  INV_X1 U454 ( .A(n588), .ZN(n585) );
  XNOR2_X2 U455 ( .A(n393), .B(KEYINPUT32), .ZN(n588) );
  XNOR2_X2 U456 ( .A(n515), .B(n514), .ZN(n600) );
  INV_X1 U457 ( .A(n630), .ZN(n636) );
  XNOR2_X2 U458 ( .A(n542), .B(n541), .ZN(n684) );
  BUF_X2 U459 ( .A(n502), .Z(n542) );
  XOR2_X1 U460 ( .A(n460), .B(KEYINPUT94), .Z(n394) );
  INV_X1 U461 ( .A(KEYINPUT64), .ZN(n628) );
  AND2_X1 U462 ( .A1(n534), .A2(n503), .ZN(n536) );
  XNOR2_X1 U463 ( .A(n752), .B(n468), .ZN(n650) );
  AND2_X1 U464 ( .A1(n640), .A2(G953), .ZN(n733) );
  XNOR2_X1 U465 ( .A(G119), .B(G110), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n395), .B(KEYINPUT95), .ZN(n401) );
  NAND2_X1 U467 ( .A1(G234), .A2(n744), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n354), .B(n397), .ZN(n430) );
  NAND2_X1 U469 ( .A1(n430), .A2(G221), .ZN(n398) );
  XNOR2_X2 U470 ( .A(G146), .B(G125), .ZN(n479) );
  XNOR2_X1 U471 ( .A(G140), .B(n750), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n731) );
  NOR2_X1 U473 ( .A1(n731), .A2(G902), .ZN(n406) );
  XOR2_X1 U474 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n404) );
  XNOR2_X1 U475 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  NAND2_X1 U476 ( .A1(n623), .A2(G234), .ZN(n402) );
  XNOR2_X1 U477 ( .A(n402), .B(KEYINPUT20), .ZN(n408) );
  NAND2_X1 U478 ( .A1(n408), .A2(G217), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U480 ( .A(n406), .B(n405), .ZN(n518) );
  AND2_X1 U481 ( .A1(n408), .A2(G221), .ZN(n410) );
  INV_X1 U482 ( .A(KEYINPUT21), .ZN(n409) );
  XNOR2_X1 U483 ( .A(n410), .B(n409), .ZN(n698) );
  NAND2_X1 U484 ( .A1(G234), .A2(G237), .ZN(n411) );
  XNOR2_X1 U485 ( .A(n411), .B(KEYINPUT14), .ZN(n681) );
  INV_X1 U486 ( .A(G902), .ZN(n458) );
  NAND2_X1 U487 ( .A1(G953), .A2(n458), .ZN(n412) );
  NAND2_X1 U488 ( .A1(n681), .A2(n412), .ZN(n509) );
  INV_X1 U489 ( .A(n509), .ZN(n415) );
  INV_X1 U490 ( .A(G952), .ZN(n640) );
  NAND2_X1 U491 ( .A1(n744), .A2(n640), .ZN(n507) );
  NAND2_X1 U492 ( .A1(G953), .A2(G900), .ZN(n413) );
  AND2_X1 U493 ( .A1(n507), .A2(n413), .ZN(n414) );
  NAND2_X1 U494 ( .A1(n415), .A2(n414), .ZN(n537) );
  NOR2_X1 U495 ( .A1(n698), .A2(n537), .ZN(n416) );
  XOR2_X1 U496 ( .A(n416), .B(KEYINPUT71), .Z(n417) );
  AND2_X1 U497 ( .A1(n407), .A2(n417), .ZN(n550) );
  INV_X1 U498 ( .A(G131), .ZN(n418) );
  XNOR2_X1 U499 ( .A(n418), .B(G140), .ZN(n460) );
  XNOR2_X1 U500 ( .A(n460), .B(n750), .ZN(n422) );
  XOR2_X1 U501 ( .A(G122), .B(G104), .Z(n420) );
  XNOR2_X1 U502 ( .A(G113), .B(G143), .ZN(n419) );
  XNOR2_X1 U503 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U504 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U505 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n424) );
  NAND2_X1 U506 ( .A1(G214), .A2(n446), .ZN(n423) );
  XNOR2_X1 U507 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U508 ( .A(n425), .B(KEYINPUT12), .Z(n426) );
  XNOR2_X1 U509 ( .A(n427), .B(n426), .ZN(n726) );
  NOR2_X1 U510 ( .A1(n726), .A2(G902), .ZN(n429) );
  XNOR2_X1 U511 ( .A(KEYINPUT13), .B(G475), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n429), .B(n428), .ZN(n544) );
  NAND2_X1 U513 ( .A1(n430), .A2(G217), .ZN(n437) );
  XNOR2_X1 U514 ( .A(G122), .B(KEYINPUT9), .ZN(n432) );
  XNOR2_X1 U515 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n431) );
  XNOR2_X1 U516 ( .A(n432), .B(n431), .ZN(n435) );
  XNOR2_X1 U517 ( .A(G116), .B(G107), .ZN(n433) );
  XNOR2_X1 U518 ( .A(n433), .B(KEYINPUT100), .ZN(n434) );
  XNOR2_X1 U519 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U520 ( .A(n437), .B(n436), .ZN(n440) );
  XNOR2_X2 U521 ( .A(KEYINPUT83), .B(G143), .ZN(n439) );
  XNOR2_X1 U522 ( .A(n440), .B(n443), .ZN(n645) );
  NAND2_X1 U523 ( .A1(n645), .A2(n458), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n441), .B(G478), .ZN(n498) );
  INV_X1 U525 ( .A(n498), .ZN(n543) );
  NAND2_X1 U526 ( .A1(n544), .A2(n543), .ZN(n669) );
  XNOR2_X1 U527 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n480) );
  XNOR2_X1 U528 ( .A(n480), .B(G137), .ZN(n442) );
  XNOR2_X1 U529 ( .A(G116), .B(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U530 ( .A(G146), .B(G131), .ZN(n448) );
  NAND2_X1 U531 ( .A1(G210), .A2(n446), .ZN(n447) );
  XNOR2_X1 U532 ( .A(n448), .B(n447), .ZN(n451) );
  XNOR2_X1 U533 ( .A(KEYINPUT66), .B(G101), .ZN(n463) );
  XNOR2_X1 U534 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n449) );
  XNOR2_X1 U535 ( .A(n463), .B(n449), .ZN(n450) );
  XNOR2_X1 U536 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U537 ( .A(n474), .B(n452), .ZN(n453) );
  XNOR2_X1 U538 ( .A(n461), .B(n453), .ZN(n637) );
  XNOR2_X2 U539 ( .A(n454), .B(G472), .ZN(n534) );
  XNOR2_X1 U540 ( .A(n534), .B(KEYINPUT6), .ZN(n599) );
  NOR2_X1 U541 ( .A1(n669), .A2(n599), .ZN(n455) );
  NAND2_X1 U542 ( .A1(n550), .A2(n455), .ZN(n456) );
  XNOR2_X1 U543 ( .A(n456), .B(KEYINPUT107), .ZN(n459) );
  INV_X1 U544 ( .A(G237), .ZN(n457) );
  NAND2_X1 U545 ( .A1(n458), .A2(n457), .ZN(n494) );
  AND2_X1 U546 ( .A1(n494), .A2(G214), .ZN(n683) );
  AND2_X1 U547 ( .A1(n459), .A2(n503), .ZN(n572) );
  XOR2_X1 U548 ( .A(G104), .B(G110), .Z(n462) );
  XNOR2_X1 U549 ( .A(n462), .B(G107), .ZN(n740) );
  XNOR2_X1 U550 ( .A(n463), .B(KEYINPUT73), .ZN(n464) );
  XNOR2_X1 U551 ( .A(n740), .B(n464), .ZN(n475) );
  XNOR2_X1 U552 ( .A(G146), .B(KEYINPUT78), .ZN(n466) );
  NAND2_X1 U553 ( .A1(n744), .A2(G227), .ZN(n465) );
  XNOR2_X1 U554 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U555 ( .A(n475), .B(n467), .ZN(n468) );
  XNOR2_X2 U556 ( .A(n469), .B(G469), .ZN(n609) );
  INV_X1 U557 ( .A(n695), .ZN(n470) );
  NAND2_X1 U558 ( .A1(n572), .A2(n470), .ZN(n471) );
  XNOR2_X1 U559 ( .A(n471), .B(KEYINPUT43), .ZN(n497) );
  XNOR2_X1 U560 ( .A(KEYINPUT16), .B(G122), .ZN(n472) );
  XNOR2_X1 U561 ( .A(n472), .B(KEYINPUT75), .ZN(n473) );
  NAND2_X1 U562 ( .A1(n744), .A2(G224), .ZN(n476) );
  XNOR2_X1 U563 ( .A(n476), .B(KEYINPUT80), .ZN(n478) );
  XNOR2_X1 U564 ( .A(KEYINPUT79), .B(KEYINPUT18), .ZN(n477) );
  XNOR2_X1 U565 ( .A(n478), .B(n477), .ZN(n484) );
  INV_X1 U566 ( .A(n484), .ZN(n482) );
  XNOR2_X1 U567 ( .A(n480), .B(n479), .ZN(n483) );
  INV_X1 U568 ( .A(n483), .ZN(n481) );
  NAND2_X1 U569 ( .A1(n482), .A2(n481), .ZN(n486) );
  NAND2_X1 U570 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U571 ( .A1(n486), .A2(n485), .ZN(n491) );
  INV_X1 U572 ( .A(n487), .ZN(n489) );
  XOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U575 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U576 ( .A1(n721), .A2(n623), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X2 U578 ( .A(n496), .B(n495), .ZN(n502) );
  NAND2_X1 U579 ( .A1(n497), .A2(n542), .ZN(n582) );
  XNOR2_X1 U580 ( .A(n582), .B(G140), .ZN(G42) );
  OR2_X1 U581 ( .A1(n544), .A2(n498), .ZN(n499) );
  XNOR2_X2 U582 ( .A(n499), .B(KEYINPUT103), .ZN(n686) );
  INV_X1 U583 ( .A(n698), .ZN(n500) );
  XNOR2_X1 U584 ( .A(n501), .B(KEYINPUT104), .ZN(n513) );
  INV_X1 U585 ( .A(n502), .ZN(n504) );
  INV_X1 U586 ( .A(n683), .ZN(n503) );
  NAND2_X1 U587 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U588 ( .A(n505), .B(KEYINPUT19), .ZN(n563) );
  NAND2_X1 U589 ( .A1(G953), .A2(G898), .ZN(n506) );
  NAND2_X1 U590 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U591 ( .A1(n509), .A2(n508), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n563), .A2(n510), .ZN(n512) );
  XNOR2_X1 U593 ( .A(KEYINPUT91), .B(KEYINPUT0), .ZN(n511) );
  XNOR2_X2 U594 ( .A(n512), .B(n511), .ZN(n525) );
  NAND2_X1 U595 ( .A1(n513), .A2(n525), .ZN(n515) );
  INV_X1 U596 ( .A(KEYINPUT22), .ZN(n514) );
  INV_X1 U597 ( .A(n534), .ZN(n608) );
  NAND2_X1 U598 ( .A1(n407), .A2(n608), .ZN(n516) );
  NOR2_X1 U599 ( .A1(n695), .A2(n516), .ZN(n517) );
  AND2_X1 U600 ( .A1(n600), .A2(n517), .ZN(n586) );
  XOR2_X1 U601 ( .A(G110), .B(n586), .Z(G12) );
  INV_X1 U602 ( .A(KEYINPUT68), .ZN(n519) );
  XNOR2_X2 U603 ( .A(n520), .B(n519), .ZN(n696) );
  INV_X1 U604 ( .A(n599), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n605), .A2(n522), .ZN(n524) );
  XNOR2_X1 U606 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n523) );
  NAND2_X1 U607 ( .A1(n682), .A2(n525), .ZN(n527) );
  XOR2_X1 U608 ( .A(KEYINPUT82), .B(KEYINPUT34), .Z(n526) );
  XNOR2_X1 U609 ( .A(n527), .B(n526), .ZN(n531) );
  INV_X1 U610 ( .A(n544), .ZN(n528) );
  OR2_X1 U611 ( .A1(n528), .A2(n543), .ZN(n561) );
  INV_X1 U612 ( .A(n561), .ZN(n529) );
  XOR2_X1 U613 ( .A(n529), .B(KEYINPUT81), .Z(n530) );
  NAND2_X1 U614 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U615 ( .A(KEYINPUT35), .ZN(n532) );
  XNOR2_X2 U616 ( .A(n533), .B(n532), .ZN(n595) );
  XNOR2_X1 U617 ( .A(n595), .B(G122), .ZN(G24) );
  XNOR2_X1 U618 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n535) );
  XNOR2_X1 U619 ( .A(n536), .B(n535), .ZN(n539) );
  INV_X1 U620 ( .A(n537), .ZN(n538) );
  AND2_X1 U621 ( .A1(n539), .A2(n356), .ZN(n540) );
  NAND2_X1 U622 ( .A1(n696), .A2(n540), .ZN(n559) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n541) );
  OR2_X1 U624 ( .A1(n544), .A2(n543), .ZN(n671) );
  OR2_X1 U625 ( .A1(n545), .A2(n671), .ZN(n581) );
  XNOR2_X1 U626 ( .A(n581), .B(G134), .ZN(G36) );
  XNOR2_X1 U627 ( .A(n557), .B(G131), .ZN(G33) );
  AND2_X1 U628 ( .A1(n695), .A2(n407), .ZN(n546) );
  AND2_X1 U629 ( .A1(n599), .A2(n546), .ZN(n547) );
  XOR2_X1 U630 ( .A(G119), .B(n585), .Z(G21) );
  INV_X1 U631 ( .A(n689), .ZN(n548) );
  NAND2_X1 U632 ( .A1(n686), .A2(n548), .ZN(n549) );
  XNOR2_X2 U633 ( .A(n549), .B(KEYINPUT41), .ZN(n714) );
  NAND2_X1 U634 ( .A1(n550), .A2(n534), .ZN(n552) );
  XOR2_X1 U635 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n551) );
  XNOR2_X1 U636 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U637 ( .A1(n553), .A2(n609), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n714), .A2(n564), .ZN(n556) );
  INV_X1 U639 ( .A(KEYINPUT111), .ZN(n554) );
  XNOR2_X1 U640 ( .A(n554), .B(KEYINPUT42), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n556), .B(n555), .ZN(n765) );
  AND2_X1 U642 ( .A1(n765), .A2(n557), .ZN(n558) );
  NOR2_X1 U643 ( .A1(n559), .A2(n542), .ZN(n560) );
  XNOR2_X1 U644 ( .A(n560), .B(KEYINPUT109), .ZN(n562) );
  OR2_X1 U645 ( .A1(n562), .A2(n561), .ZN(n664) );
  AND2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n666) );
  AND2_X1 U647 ( .A1(n669), .A2(n671), .ZN(n688) );
  INV_X1 U648 ( .A(n688), .ZN(n613) );
  NAND2_X1 U649 ( .A1(n666), .A2(n613), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n565), .A2(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U651 ( .A1(n664), .A2(n566), .ZN(n568) );
  INV_X1 U652 ( .A(KEYINPUT84), .ZN(n567) );
  XNOR2_X1 U653 ( .A(n568), .B(n567), .ZN(n579) );
  NOR2_X1 U654 ( .A1(KEYINPUT47), .A2(n688), .ZN(n569) );
  XNOR2_X1 U655 ( .A(n569), .B(KEYINPUT76), .ZN(n570) );
  NAND2_X1 U656 ( .A1(n666), .A2(n570), .ZN(n577) );
  INV_X1 U657 ( .A(n542), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U659 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n575), .A2(n695), .ZN(n576) );
  XNOR2_X1 U662 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n580) );
  AND2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U664 ( .A1(n753), .A2(n623), .ZN(n622) );
  INV_X1 U665 ( .A(KEYINPUT67), .ZN(n584) );
  INV_X1 U666 ( .A(n586), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n590) );
  INV_X1 U668 ( .A(KEYINPUT88), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n590), .B(n589), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n591), .A2(n594), .ZN(n593) );
  INV_X1 U671 ( .A(KEYINPUT44), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n593), .B(n592), .ZN(n620) );
  INV_X1 U673 ( .A(n594), .ZN(n598) );
  INV_X1 U674 ( .A(n595), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n596), .A2(KEYINPUT67), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n618) );
  AND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n695), .A2(n407), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U680 ( .A(KEYINPUT105), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n604), .B(n603), .ZN(n762) );
  AND2_X1 U682 ( .A1(n605), .A2(n534), .ZN(n704) );
  NAND2_X1 U683 ( .A1(n704), .A2(n525), .ZN(n607) );
  XNOR2_X1 U684 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n607), .B(n606), .ZN(n668) );
  NAND2_X1 U686 ( .A1(n696), .A2(n608), .ZN(n611) );
  INV_X1 U687 ( .A(n609), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U689 ( .A1(n612), .A2(n525), .ZN(n655) );
  OR2_X1 U690 ( .A1(n668), .A2(n655), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT102), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n762), .A2(n616), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT45), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n622), .A2(n631), .ZN(n627) );
  INV_X1 U698 ( .A(n623), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n624), .A2(KEYINPUT2), .ZN(n625) );
  XOR2_X1 U700 ( .A(KEYINPUT65), .B(n625), .Z(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n630) );
  INV_X1 U703 ( .A(n734), .ZN(n634) );
  INV_X1 U704 ( .A(n753), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n632), .A2(KEYINPUT2), .ZN(n633) );
  NOR2_X2 U706 ( .A1(n634), .A2(n633), .ZN(n679) );
  INV_X1 U707 ( .A(n679), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n725), .A2(G472), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n637), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n641) );
  XNOR2_X1 U711 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(G57) );
  NAND2_X1 U713 ( .A1(n729), .A2(G478), .ZN(n644) );
  XOR2_X1 U714 ( .A(n645), .B(n644), .Z(n646) );
  NOR2_X1 U715 ( .A1(n646), .A2(n733), .ZN(G63) );
  NAND2_X1 U716 ( .A1(n725), .A2(G469), .ZN(n652) );
  XNOR2_X1 U717 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n648) );
  XNOR2_X1 U718 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT120), .ZN(G54) );
  INV_X1 U723 ( .A(n655), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n657), .A2(n669), .ZN(n656) );
  XOR2_X1 U725 ( .A(G104), .B(n656), .Z(G6) );
  NOR2_X1 U726 ( .A1(n657), .A2(n671), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(G107), .B(n660), .ZN(G9) );
  XOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .Z(n663) );
  INV_X1 U731 ( .A(n671), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n666), .A2(n661), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G30) );
  XNOR2_X1 U734 ( .A(G143), .B(KEYINPUT114), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(G45) );
  NAND2_X1 U736 ( .A1(n666), .A2(n372), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(G146), .ZN(G48) );
  INV_X1 U738 ( .A(n668), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n672), .A2(n669), .ZN(n670) );
  XOR2_X1 U740 ( .A(G113), .B(n670), .Z(G15) );
  NOR2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U742 ( .A(G116), .B(n673), .Z(G18) );
  OR2_X1 U743 ( .A1(n734), .A2(KEYINPUT2), .ZN(n677) );
  INV_X1 U744 ( .A(KEYINPUT2), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n753), .A2(n674), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT86), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n680), .A2(G953), .ZN(n719) );
  NAND2_X1 U750 ( .A1(G952), .A2(n681), .ZN(n713) );
  INV_X1 U751 ( .A(n715), .ZN(n693) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U754 ( .A(KEYINPUT116), .B(n687), .Z(n691) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U758 ( .A(n694), .B(KEYINPUT117), .ZN(n710) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U760 ( .A(KEYINPUT50), .B(n697), .Z(n703) );
  XOR2_X1 U761 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n700) );
  NAND2_X1 U762 ( .A1(n698), .A2(n407), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n701), .A2(n534), .ZN(n702) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n706) );
  INV_X1 U766 ( .A(n704), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U768 ( .A(KEYINPUT51), .B(n707), .Z(n708) );
  NAND2_X1 U769 ( .A1(n708), .A2(n714), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT52), .B(n711), .Z(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n717) );
  AND2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U776 ( .A(KEYINPUT53), .B(n720), .Z(G75) );
  XNOR2_X1 U777 ( .A(KEYINPUT55), .B(KEYINPUT90), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT54), .ZN(n723) );
  XNOR2_X1 U779 ( .A(n721), .B(n723), .ZN(n724) );
  XNOR2_X1 U780 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT93), .ZN(n727) );
  NAND2_X1 U782 ( .A1(n729), .A2(G217), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(G66) );
  NAND2_X1 U785 ( .A1(n734), .A2(n744), .ZN(n739) );
  NAND2_X1 U786 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n735), .B(KEYINPUT61), .ZN(n736) );
  XNOR2_X1 U788 ( .A(KEYINPUT122), .B(n736), .ZN(n737) );
  NAND2_X1 U789 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n749) );
  XOR2_X1 U791 ( .A(n740), .B(KEYINPUT123), .Z(n742) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n743), .B(G101), .ZN(n746) );
  NOR2_X1 U794 ( .A1(n744), .A2(G898), .ZN(n745) );
  NOR2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U796 ( .A(KEYINPUT124), .B(n747), .ZN(n748) );
  XNOR2_X1 U797 ( .A(n749), .B(n748), .ZN(G69) );
  XOR2_X1 U798 ( .A(KEYINPUT125), .B(n750), .Z(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(n755) );
  XOR2_X1 U800 ( .A(n755), .B(n753), .Z(n754) );
  NOR2_X1 U801 ( .A1(n754), .A2(G953), .ZN(n760) );
  XNOR2_X1 U802 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U804 ( .A1(G953), .A2(n757), .ZN(n758) );
  XOR2_X1 U805 ( .A(KEYINPUT126), .B(n758), .Z(n759) );
  NOR2_X1 U806 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U807 ( .A(KEYINPUT127), .B(n761), .ZN(G72) );
  XNOR2_X1 U808 ( .A(G101), .B(n762), .ZN(G3) );
  XOR2_X1 U809 ( .A(G125), .B(n763), .Z(n764) );
  XNOR2_X1 U810 ( .A(KEYINPUT37), .B(n764), .ZN(G27) );
  XNOR2_X1 U811 ( .A(G137), .B(n765), .ZN(G39) );
endmodule

