//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n190), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(G146), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G110), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(KEYINPUT24), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT24), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT74), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT24), .B(G110), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT75), .ZN(new_n209));
  OAI211_X1 g023(.A(G119), .B(new_n206), .C1(new_n209), .C2(KEYINPUT23), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n204), .B2(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT75), .B1(new_n204), .B2(G128), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n196), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n203), .A2(new_n208), .B1(KEYINPUT76), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n196), .A4(new_n210), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n195), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n208), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n199), .A2(new_n202), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G110), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n224));
  AOI21_X1  g038(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n221), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT77), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n203), .A2(new_n208), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(KEYINPUT76), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n218), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n195), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n226), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT22), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(G137), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n226), .A3(new_n239), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT25), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n241), .A2(new_n246), .A3(new_n242), .A4(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(G217), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(G234), .B2(new_n242), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n241), .A2(new_n243), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n249), .A2(G902), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT26), .B(G101), .Z(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G137), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n262), .C2(G137), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G134), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT11), .B1(new_n270), .B2(KEYINPUT65), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n269), .A2(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(new_n262), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n273), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n277), .B2(new_n264), .ZN(new_n278));
  INV_X1    g092(.A(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G143), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G128), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT64), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n286), .ZN(new_n290));
  NOR2_X1   g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G143), .B(G146), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(KEYINPUT64), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n278), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n265), .B1(new_n276), .B2(new_n267), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n264), .B1(new_n270), .B2(new_n263), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n280), .A3(new_n282), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n281), .A2(KEYINPUT1), .A3(G146), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n300), .B(new_n301), .C1(G128), .C2(new_n293), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT66), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  AND4_X1   g118(.A1(KEYINPUT66), .A2(new_n272), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n295), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G119), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n204), .A2(KEYINPUT67), .A3(G116), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n309), .A2(new_n310), .B1(new_n308), .B2(G119), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT2), .A2(G113), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT2), .A2(G113), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(G119), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n316), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n306), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n285), .A2(new_n287), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n278), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT68), .B1(new_n315), .B2(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n317), .ZN(new_n325));
  INV_X1    g139(.A(new_n314), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n311), .A2(new_n314), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n272), .A2(new_n302), .A3(new_n304), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n323), .A2(new_n324), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n261), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n260), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n323), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n272), .A2(new_n302), .A3(KEYINPUT66), .A4(new_n304), .ZN(new_n341));
  INV_X1    g155(.A(new_n294), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(new_n288), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n340), .A2(new_n341), .B1(new_n343), .B2(new_n278), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n320), .B(new_n338), .C1(new_n344), .C2(KEYINPUT30), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n263), .B1(new_n268), .B2(new_n271), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n296), .B1(new_n346), .B2(G131), .ZN(new_n347));
  INV_X1    g161(.A(new_n322), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n331), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n324), .A2(new_n330), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n260), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT31), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n337), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(G472), .A2(G902), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n358), .B(KEYINPUT71), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT32), .B1(new_n357), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n260), .B1(new_n332), .B2(new_n334), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n333), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n260), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n345), .B2(new_n332), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n364), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n261), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n340), .A2(new_n341), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n319), .B1(new_n373), .B2(new_n295), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n374), .B2(new_n351), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n375), .B2(new_n366), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n345), .A2(new_n332), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n260), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT72), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n349), .A2(new_n350), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n334), .B1(new_n380), .B2(new_n332), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(KEYINPUT73), .A3(KEYINPUT29), .A4(new_n366), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT73), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n335), .A2(KEYINPUT29), .A3(new_n369), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n371), .A2(new_n379), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G472), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n254), .B1(new_n363), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT78), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G221), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT79), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G140), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n236), .A2(G227), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT80), .A3(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(new_n401), .A3(KEYINPUT80), .A4(G104), .ZN(new_n405));
  INV_X1    g219(.A(G104), .ZN(new_n406));
  AOI21_X1  g220(.A(G101), .B1(new_n406), .B2(G107), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n406), .A2(G107), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n401), .A2(G104), .ZN(new_n410));
  OAI21_X1  g224(.A(G101), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n400), .B1(new_n412), .B2(new_n302), .ZN(new_n413));
  AND4_X1   g227(.A1(new_n400), .A2(new_n302), .A3(new_n408), .A4(new_n411), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n413), .A2(new_n414), .B1(new_n302), .B2(new_n412), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT12), .A3(new_n278), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n302), .B1(new_n408), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n301), .B1(new_n293), .B2(G128), .ZN(new_n419));
  INV_X1    g233(.A(new_n300), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n408), .A2(new_n411), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT81), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n302), .A2(new_n400), .A3(new_n408), .A4(new_n411), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n417), .B1(new_n425), .B2(new_n347), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n410), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n403), .A2(new_n405), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G101), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT4), .A3(G101), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n421), .A2(new_n422), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n434), .A2(new_n322), .B1(KEYINPUT10), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n413), .B2(new_n414), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n438), .A3(new_n347), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n399), .B1(new_n427), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(KEYINPUT4), .A2(new_n408), .B1(new_n429), .B2(G101), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n429), .A2(KEYINPUT4), .A3(G101), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n322), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT10), .B1(new_n423), .B2(new_n424), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n278), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n439), .A3(new_n399), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT82), .B1(new_n440), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT12), .B1(new_n415), .B2(new_n278), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n425), .A2(new_n417), .A3(new_n347), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n439), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n398), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n448), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n456), .A3(G469), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n242), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n447), .A2(new_n439), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n398), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n439), .B(new_n399), .C1(new_n451), .C2(new_n452), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n395), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G475), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n256), .A2(G214), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT88), .A3(G143), .ZN(new_n468));
  OR2_X1    g282(.A1(KEYINPUT88), .A2(G143), .ZN(new_n469));
  NAND2_X1  g283(.A1(KEYINPUT88), .A2(G143), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(G214), .A3(new_n256), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(KEYINPUT18), .A2(G131), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n194), .A2(G146), .ZN(new_n475));
  XNOR2_X1  g289(.A(G125), .B(G140), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n279), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n472), .A2(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n473), .B1(new_n468), .B2(new_n471), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n468), .A2(new_n471), .A3(KEYINPUT17), .A4(G131), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n191), .A2(new_n192), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n279), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n483), .A3(new_n193), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n472), .A2(new_n264), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n468), .A2(G131), .A3(new_n471), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n486), .A4(new_n487), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n480), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G113), .B(G122), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n406), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n466), .B1(new_n495), .B2(new_n242), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n468), .A2(G131), .A3(new_n471), .ZN(new_n498));
  AOI21_X1  g312(.A(G131), .B1(new_n468), .B2(new_n471), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n485), .A2(KEYINPUT89), .A3(new_n487), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT19), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n194), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n476), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n224), .B1(new_n506), .B2(new_n279), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n478), .A2(new_n479), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n494), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n494), .B1(new_n508), .B2(new_n509), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n488), .A2(new_n489), .ZN(new_n517));
  INV_X1    g331(.A(new_n484), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n491), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n494), .A3(new_n509), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT93), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(KEYINPUT91), .B2(new_n515), .ZN(new_n529));
  INV_X1    g343(.A(new_n516), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(new_n523), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n496), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G214), .B1(G237), .B2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G210), .B1(G237), .B2(G902), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n283), .A2(new_n206), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n538), .A2(new_n189), .A3(new_n300), .A4(new_n301), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n285), .A2(G125), .A3(new_n287), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n537), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G224), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n543), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n434), .A2(new_n320), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT5), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n204), .A3(G116), .ZN(new_n549));
  OAI211_X1 g363(.A(G113), .B(new_n549), .C1(new_n325), .C2(new_n548), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n412), .A3(new_n329), .ZN(new_n551));
  XOR2_X1   g365(.A(G110), .B(G122), .Z(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT83), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n551), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT84), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(KEYINPUT6), .A3(new_n558), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n546), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n545), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT7), .B(new_n563), .C1(new_n543), .C2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n553), .B(KEYINPUT8), .ZN(new_n566));
  INV_X1    g380(.A(new_n551), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n412), .B1(new_n550), .B2(new_n329), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(KEYINPUT7), .ZN(new_n570));
  OAI221_X1 g384(.A(new_n570), .B1(KEYINPUT86), .B2(new_n545), .C1(new_n541), .C2(new_n542), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n565), .A2(new_n569), .A3(new_n554), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n242), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n536), .B1(new_n562), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  INV_X1    g389(.A(new_n546), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n554), .A2(KEYINPUT6), .B1(new_n556), .B2(new_n558), .ZN(new_n577));
  INV_X1    g391(.A(new_n561), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n579), .A3(new_n535), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n534), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT15), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n236), .A2(G217), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n392), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G128), .B(G143), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT13), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n281), .A2(G128), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n586), .B(G134), .C1(KEYINPUT13), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(G116), .B(G122), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n401), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n262), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n585), .B(new_n262), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n308), .A2(KEYINPUT14), .A3(G122), .ZN(new_n594));
  INV_X1    g408(.A(new_n589), .ZN(new_n595));
  OAI211_X1 g409(.A(G107), .B(new_n594), .C1(new_n595), .C2(KEYINPUT14), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n589), .A2(new_n401), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n584), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n592), .A2(new_n598), .A3(new_n584), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT94), .B1(new_n602), .B2(new_n242), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  OAI211_X1 g418(.A(KEYINPUT94), .B(new_n242), .C1(new_n604), .C2(new_n599), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n582), .B(G478), .C1(new_n603), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n582), .A2(G478), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n242), .B(new_n608), .C1(new_n604), .C2(new_n599), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT95), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G952), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n612), .A2(KEYINPUT96), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(KEYINPUT96), .ZN(new_n614));
  AOI21_X1  g428(.A(G953), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT21), .B(G898), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n532), .A2(new_n581), .A3(new_n611), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n390), .A2(new_n465), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NOR2_X1   g438(.A1(new_n604), .A2(new_n599), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT97), .B1(new_n592), .B2(new_n598), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  OAI22_X1  g443(.A1(new_n604), .A2(new_n599), .B1(new_n626), .B2(new_n627), .ZN(new_n630));
  AND4_X1   g444(.A1(G478), .A2(new_n629), .A3(new_n242), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n625), .B2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(G478), .B1(new_n633), .B2(new_n605), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n523), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n512), .A2(new_n513), .B1(new_n492), .B2(new_n494), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n516), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n531), .B1(new_n638), .B2(new_n525), .ZN(new_n639));
  INV_X1    g453(.A(new_n496), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n581), .A2(new_n621), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n369), .B1(new_n375), .B2(new_n335), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n345), .A2(new_n355), .A3(new_n352), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n355), .B1(new_n345), .B2(new_n352), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n359), .ZN(new_n649));
  INV_X1    g463(.A(G472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n357), .B2(new_n242), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n649), .A2(new_n651), .A3(new_n254), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n644), .A2(new_n465), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  NOR2_X1   g469(.A1(new_n611), .A2(new_n496), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n638), .A2(new_n525), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n527), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n638), .A2(KEYINPUT98), .A3(new_n525), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n643), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n465), .A3(new_n652), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT99), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n651), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  INV_X1    g482(.A(new_n252), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n219), .A2(new_n227), .A3(KEYINPUT77), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n234), .B1(new_n233), .B2(new_n226), .ZN(new_n671));
  OAI22_X1  g485(.A1(new_n670), .A2(new_n671), .B1(KEYINPUT36), .B2(new_n240), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n240), .A2(KEYINPUT36), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n228), .A2(new_n235), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n249), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n244), .B2(KEYINPUT25), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n668), .B(new_n675), .C1(new_n677), .C2(new_n247), .ZN(new_n678));
  INV_X1    g492(.A(new_n675), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n250), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n622), .A2(new_n465), .A3(new_n667), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  AND2_X1   g498(.A1(new_n681), .A2(new_n465), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n574), .A2(new_n580), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n533), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n363), .B2(new_n389), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n617), .B(KEYINPUT102), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n620), .A2(G900), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n656), .A2(new_n659), .A3(new_n660), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n685), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  OR2_X1    g510(.A1(new_n686), .A2(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(KEYINPUT103), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT32), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n648), .B2(new_n359), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n360), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n260), .B1(new_n345), .B2(new_n332), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n380), .A2(new_n332), .A3(new_n260), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n242), .ZN(new_n707));
  OAI21_X1  g521(.A(G472), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n703), .A2(KEYINPUT104), .A3(new_n704), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n697), .A2(KEYINPUT38), .A3(new_n698), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n675), .B1(new_n677), .B2(new_n247), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n532), .A2(new_n716), .A3(new_n611), .A4(new_n534), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n701), .A2(new_n713), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n692), .B(KEYINPUT105), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT39), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n465), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT40), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n718), .B2(new_n722), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n281), .ZN(G45));
  INV_X1    g541(.A(new_n692), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n532), .A2(new_n635), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n685), .A2(new_n688), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NOR2_X1   g545(.A1(new_n445), .A2(new_n446), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n398), .B1(new_n732), .B2(new_n347), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n427), .A2(new_n733), .B1(new_n460), .B2(new_n398), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n734), .B2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n461), .A2(new_n462), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n458), .A3(new_n242), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n735), .A2(new_n394), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n390), .A2(new_n644), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n390), .A2(new_n662), .A3(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  AND2_X1   g557(.A1(new_n738), .A2(new_n621), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n532), .A3(new_n611), .A4(new_n681), .ZN(new_n745));
  INV_X1    g559(.A(new_n688), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n204), .ZN(G21));
  NOR3_X1   g562(.A1(new_n687), .A2(new_n532), .A3(new_n611), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n646), .A2(new_n647), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n260), .B1(new_n336), .B2(new_n381), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n359), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n651), .A2(new_n254), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n744), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT107), .Z(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n738), .A2(new_n581), .A3(new_n641), .A4(new_n692), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n651), .A2(new_n715), .A3(new_n752), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n735), .A2(new_n394), .A3(new_n737), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n687), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n651), .A2(new_n752), .A3(new_n715), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n729), .A3(KEYINPUT108), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  AOI22_X1  g580(.A1(new_n416), .A2(new_n426), .B1(new_n732), .B2(new_n347), .ZN(new_n767));
  OAI211_X1 g581(.A(G469), .B(new_n448), .C1(new_n767), .C2(new_n399), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n454), .A2(KEYINPUT110), .A3(G469), .A4(new_n448), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n459), .B(KEYINPUT109), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n737), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n772), .B1(new_n463), .B2(new_n458), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n771), .A4(new_n770), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n775), .A2(new_n394), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n686), .A2(new_n534), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n390), .A3(new_n729), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  INV_X1    g598(.A(new_n254), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n388), .A2(G472), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n703), .A2(new_n704), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n785), .B(new_n780), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT42), .A3(new_n729), .A4(new_n779), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n784), .B1(new_n783), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G131), .ZN(G33));
  NAND3_X1  g608(.A1(new_n775), .A2(new_n394), .A3(new_n778), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n788), .A2(new_n795), .A3(new_n693), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n262), .ZN(G36));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n450), .B2(new_n456), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n454), .A2(KEYINPUT45), .A3(new_n448), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(G469), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n802), .B2(new_n772), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT46), .B(new_n773), .C1(new_n799), .C2(new_n801), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n737), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n394), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT113), .B1(new_n807), .B2(new_n720), .ZN(new_n808));
  AND4_X1   g622(.A1(KEYINPUT113), .A2(new_n805), .A3(new_n394), .A4(new_n720), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n532), .B1(new_n634), .B2(new_n631), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT43), .Z(new_n812));
  INV_X1    g626(.A(new_n667), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n716), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(KEYINPUT44), .A3(new_n813), .A4(new_n716), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n780), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n269), .ZN(G39));
  OR2_X1    g634(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n389), .A2(new_n703), .A3(new_n704), .ZN(new_n823));
  INV_X1    g637(.A(new_n780), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n785), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n729), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND2_X1  g641(.A1(new_n701), .A2(new_n714), .ZN(new_n828));
  INV_X1    g642(.A(new_n713), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n735), .A2(new_n737), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT49), .Z(new_n831));
  NOR4_X1   g645(.A1(new_n811), .A2(new_n254), .A3(new_n395), .A4(new_n534), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT114), .Z(new_n834));
  INV_X1    g648(.A(new_n689), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n812), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n753), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n533), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n828), .A2(new_n738), .A3(new_n841), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n837), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n824), .A2(new_n761), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n763), .A3(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n824), .A2(new_n254), .A3(new_n761), .A4(new_n617), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n829), .A2(new_n847), .A3(new_n532), .A4(new_n635), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n843), .A2(new_n844), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n836), .A2(new_n753), .A3(new_n780), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n821), .A2(new_n822), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n735), .A2(new_n395), .A3(new_n737), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n836), .A2(new_n390), .A3(new_n845), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT48), .Z(new_n860));
  NAND3_X1  g674(.A1(new_n829), .A2(new_n641), .A3(new_n847), .ZN(new_n861));
  INV_X1    g675(.A(new_n762), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n615), .B(new_n861), .C1(new_n837), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n855), .B(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n849), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n858), .B(new_n864), .C1(KEYINPUT51), .C2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n739), .A2(new_n742), .A3(new_n623), .A4(new_n682), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n607), .A2(new_n610), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n532), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n642), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n643), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n465), .A4(new_n652), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n754), .B(new_n874), .C1(new_n745), .C2(new_n746), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n791), .A3(new_n792), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n639), .A2(new_n640), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n250), .A2(new_n880), .A3(new_n679), .A4(new_n692), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n581), .A2(new_n879), .A3(new_n881), .A4(new_n870), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n715), .B2(new_n692), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n713), .A2(new_n779), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n685), .B(new_n688), .C1(new_n694), .C2(new_n729), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n765), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n765), .A2(new_n885), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n870), .A2(new_n496), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n659), .A2(new_n660), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n823), .A2(new_n893), .A3(new_n465), .A4(new_n681), .ZN(new_n894));
  INV_X1    g708(.A(new_n394), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n774), .B2(KEYINPUT111), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n641), .A3(new_n763), .A4(new_n778), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n780), .A2(new_n692), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n789), .A2(new_n694), .A3(new_n779), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n894), .B2(new_n897), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n904), .A2(new_n796), .A3(KEYINPUT115), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n888), .B(new_n890), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n878), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n783), .A2(new_n790), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n876), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n912), .B2(new_n906), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n888), .A2(new_n890), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n891), .A3(new_n902), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT115), .B1(new_n904), .B2(new_n796), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n913), .B1(new_n783), .B2(new_n790), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n917), .A2(new_n920), .A3(new_n876), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n868), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n834), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n236), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n921), .A2(new_n876), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n906), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n793), .A2(new_n917), .A3(new_n920), .A4(new_n876), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n913), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n242), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n577), .A2(new_n578), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n546), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n579), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  OAI21_X1  g754(.A(new_n930), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT120), .B1(new_n934), .B2(new_n242), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n916), .A2(new_n922), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(G902), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n535), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT121), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n943), .B2(G902), .ZN(new_n950));
  AOI211_X1 g764(.A(KEYINPUT120), .B(new_n242), .C1(new_n916), .C2(new_n922), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n536), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n953), .A3(new_n947), .A4(new_n940), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n941), .B1(new_n949), .B2(new_n954), .ZN(G51));
  NAND2_X1  g769(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n924), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n772), .B(KEYINPUT57), .Z(new_n959));
  OAI21_X1  g773(.A(new_n736), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n802), .B1(new_n950), .B2(new_n951), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n929), .B1(new_n960), .B2(new_n961), .ZN(G54));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n950), .B2(new_n951), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n516), .A3(new_n637), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n521), .B(new_n963), .C1(new_n950), .C2(new_n951), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n965), .A2(new_n930), .A3(new_n966), .ZN(G60));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n629), .A2(new_n630), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT59), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n925), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n969), .A2(new_n971), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n916), .A2(new_n923), .A3(new_n922), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n923), .B1(new_n916), .B2(new_n922), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n930), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n968), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n907), .A2(new_n878), .A3(KEYINPUT53), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n923), .B1(new_n979), .B2(new_n916), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n971), .B1(new_n980), .B2(new_n974), .ZN(new_n981));
  INV_X1    g795(.A(new_n969), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(KEYINPUT122), .A3(new_n930), .A4(new_n976), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n978), .A2(new_n984), .ZN(G63));
  INV_X1    g799(.A(new_n672), .ZN(new_n986));
  INV_X1    g800(.A(new_n674), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  OR3_X1    g804(.A1(new_n934), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n934), .A2(new_n990), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n991), .B(new_n930), .C1(new_n251), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n992), .A2(new_n251), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n991), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(G66));
  NAND2_X1  g812(.A1(new_n877), .A2(new_n236), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  OAI21_X1  g814(.A(G953), .B1(new_n618), .B2(new_n544), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n937), .B1(G898), .B2(new_n236), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  OAI21_X1  g819(.A(new_n338), .B1(new_n344), .B2(KEYINPUT30), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n506), .B(KEYINPUT125), .Z(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G900), .A2(G953), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n810), .A2(new_n818), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n765), .A2(new_n886), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n826), .A2(new_n902), .A3(new_n1011), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n390), .B(new_n749), .C1(new_n808), .C2(new_n809), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1010), .A2(new_n1012), .A3(new_n793), .A4(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1008), .B(new_n1009), .C1(new_n1014), .C2(G953), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n721), .B(new_n788), .C1(new_n642), .C2(new_n871), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n826), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT62), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n724), .A2(new_n1020), .A3(new_n725), .A4(new_n1011), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n724), .A2(new_n725), .A3(new_n1011), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1010), .A2(new_n1019), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n819), .A2(new_n1018), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1027), .A2(KEYINPUT126), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1028));
  AOI21_X1  g842(.A(G953), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1015), .B1(new_n1029), .B2(new_n1008), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n236), .B1(G227), .B2(G900), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1031), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1033), .B(new_n1015), .C1(new_n1029), .C2(new_n1008), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1034), .ZN(G72));
  XNOR2_X1  g849(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n650), .A2(new_n242), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1039), .B1(new_n1014), .B2(new_n877), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n377), .A2(new_n369), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n1041), .A2(new_n705), .A3(new_n1038), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1043), .B1(new_n908), .B2(new_n914), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1042), .A2(new_n930), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1026), .A2(new_n1028), .A3(new_n876), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n1039), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1045), .B1(new_n705), .B2(new_n1047), .ZN(G57));
endmodule


