

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751;

  NOR2_X1 U368 ( .A1(n634), .A2(n720), .ZN(n408) );
  NOR2_X1 U369 ( .A1(n705), .A2(n720), .ZN(n409) );
  NOR2_X1 U370 ( .A1(n627), .A2(n720), .ZN(n629) );
  XNOR2_X1 U371 ( .A(n714), .B(n715), .ZN(n347) );
  INV_X1 U372 ( .A(KEYINPUT102), .ZN(n351) );
  XNOR2_X1 U373 ( .A(n396), .B(KEYINPUT31), .ZN(n657) );
  NOR2_X1 U374 ( .A1(n347), .A2(n720), .ZN(G63) );
  XNOR2_X2 U375 ( .A(n348), .B(n473), .ZN(n373) );
  XNOR2_X2 U376 ( .A(n527), .B(n447), .ZN(n348) );
  NAND2_X1 U377 ( .A1(n350), .A2(n349), .ZN(n544) );
  INV_X1 U378 ( .A(n636), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n542), .B(n351), .ZN(n350) );
  INV_X1 U380 ( .A(G953), .ZN(n743) );
  NOR2_X2 U381 ( .A1(n675), .A2(n590), .ZN(n612) );
  NOR2_X1 U382 ( .A1(n539), .A2(n538), .ZN(n656) );
  NOR2_X2 U383 ( .A1(n377), .A2(n748), .ZN(n364) );
  XNOR2_X1 U384 ( .A(n395), .B(n394), .ZN(n696) );
  XNOR2_X2 U385 ( .A(n433), .B(n461), .ZN(n562) );
  NOR2_X2 U386 ( .A1(n546), .A2(KEYINPUT44), .ZN(n554) );
  XNOR2_X2 U387 ( .A(n373), .B(n517), .ZN(n482) );
  NOR2_X1 U388 ( .A1(n429), .A2(n427), .ZN(n426) );
  NOR2_X1 U389 ( .A1(n696), .A2(n430), .ZN(n429) );
  XNOR2_X1 U390 ( .A(n607), .B(KEYINPUT82), .ZN(n602) );
  NOR2_X2 U391 ( .A1(n680), .A2(n679), .ZN(n540) );
  XNOR2_X1 U392 ( .A(n480), .B(n479), .ZN(n563) );
  XNOR2_X1 U393 ( .A(n728), .B(n380), .ZN(n702) );
  AND2_X1 U394 ( .A1(n422), .A2(n437), .ZN(n710) );
  AND2_X1 U395 ( .A1(n437), .A2(G475), .ZN(n413) );
  AND2_X1 U396 ( .A1(n437), .A2(G210), .ZN(n414) );
  AND2_X1 U397 ( .A1(n437), .A2(G472), .ZN(n412) );
  XNOR2_X1 U398 ( .A(n472), .B(KEYINPUT0), .ZN(n431) );
  NOR2_X1 U399 ( .A1(n597), .A2(n471), .ZN(n472) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n523) );
  XNOR2_X1 U401 ( .A(n415), .B(G125), .ZN(n501) );
  INV_X1 U402 ( .A(G146), .ZN(n415) );
  INV_X1 U403 ( .A(n663), .ZN(n619) );
  XNOR2_X1 U404 ( .A(n370), .B(n611), .ZN(n621) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n611) );
  AND2_X1 U406 ( .A1(n606), .A2(n391), .ZN(n370) );
  XNOR2_X1 U407 ( .A(n577), .B(n493), .ZN(n680) );
  INV_X1 U408 ( .A(KEYINPUT1), .ZN(n493) );
  NOR2_X1 U409 ( .A1(n624), .A2(G902), .ZN(n480) );
  XOR2_X1 U410 ( .A(KEYINPUT16), .B(KEYINPUT75), .Z(n450) );
  XNOR2_X1 U411 ( .A(n444), .B(KEYINPUT22), .ZN(n550) );
  INV_X1 U412 ( .A(n675), .ZN(n445) );
  INV_X1 U413 ( .A(n602), .ZN(n601) );
  XOR2_X1 U414 ( .A(KEYINPUT69), .B(G137), .Z(n473) );
  XNOR2_X1 U415 ( .A(G119), .B(G146), .ZN(n475) );
  XNOR2_X1 U416 ( .A(n452), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U417 ( .A(n355), .B(n451), .ZN(n452) );
  XNOR2_X1 U418 ( .A(G113), .B(G101), .ZN(n451) );
  NAND2_X1 U419 ( .A1(G234), .A2(n743), .ZN(n505) );
  XNOR2_X1 U420 ( .A(n443), .B(G122), .ZN(n521) );
  INV_X1 U421 ( .A(G104), .ZN(n443) );
  XNOR2_X1 U422 ( .A(G143), .B(G113), .ZN(n522) );
  XOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  XNOR2_X1 U424 ( .A(n483), .B(n457), .ZN(n382) );
  XNOR2_X1 U425 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n454) );
  XOR2_X1 U426 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n455) );
  NAND2_X1 U427 ( .A1(n369), .A2(n368), .ZN(n742) );
  INV_X1 U428 ( .A(n620), .ZN(n368) );
  INV_X1 U429 ( .A(KEYINPUT45), .ZN(n560) );
  XOR2_X1 U430 ( .A(KEYINPUT73), .B(KEYINPUT24), .Z(n507) );
  XNOR2_X1 U431 ( .A(G128), .B(KEYINPUT94), .ZN(n506) );
  XNOR2_X1 U432 ( .A(n500), .B(KEYINPUT23), .ZN(n504) );
  XNOR2_X1 U433 ( .A(n503), .B(n502), .ZN(n735) );
  XOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n502) );
  BUF_X1 U435 ( .A(n696), .Z(n400) );
  XNOR2_X1 U436 ( .A(n460), .B(KEYINPUT79), .ZN(n461) );
  NAND2_X1 U437 ( .A1(n702), .A2(n622), .ZN(n433) );
  NOR2_X1 U438 ( .A1(n667), .A2(n668), .ZN(n579) );
  XNOR2_X1 U439 ( .A(n573), .B(n572), .ZN(n617) );
  XNOR2_X1 U440 ( .A(n571), .B(KEYINPUT84), .ZN(n572) );
  AND2_X1 U441 ( .A1(n665), .A2(n584), .ZN(n573) );
  XNOR2_X1 U442 ( .A(n481), .B(KEYINPUT6), .ZN(n589) );
  XNOR2_X1 U443 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U444 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n418) );
  OR2_X1 U445 ( .A1(n405), .A2(KEYINPUT104), .ZN(n385) );
  INV_X1 U446 ( .A(n416), .ZN(n398) );
  AND2_X1 U447 ( .A1(n577), .A2(n407), .ZN(n570) );
  INV_X1 U448 ( .A(n679), .ZN(n407) );
  OR2_X1 U449 ( .A1(n718), .A2(G902), .ZN(n411) );
  INV_X1 U450 ( .A(KEYINPUT4), .ZN(n447) );
  AND2_X1 U451 ( .A1(n546), .A2(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U452 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n410) );
  XNOR2_X1 U453 ( .A(n442), .B(G110), .ZN(n499) );
  INV_X1 U454 ( .A(G119), .ZN(n442) );
  XNOR2_X1 U455 ( .A(G146), .B(G110), .ZN(n484) );
  XNOR2_X1 U456 ( .A(n482), .B(KEYINPUT93), .ZN(n734) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .ZN(n622) );
  NOR2_X1 U458 ( .A1(G902), .A2(G237), .ZN(n459) );
  XNOR2_X1 U459 ( .A(KEYINPUT38), .B(n586), .ZN(n665) );
  NOR2_X1 U460 ( .A1(n392), .A2(n675), .ZN(n575) );
  AND2_X1 U461 ( .A1(n405), .A2(KEYINPUT104), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n482), .B(n371), .ZN(n624) );
  XNOR2_X1 U463 ( .A(n478), .B(n372), .ZN(n371) );
  XNOR2_X1 U464 ( .A(n477), .B(n352), .ZN(n372) );
  XNOR2_X1 U465 ( .A(n474), .B(G134), .ZN(n517) );
  XNOR2_X1 U466 ( .A(n528), .B(n402), .ZN(n630) );
  XNOR2_X1 U467 ( .A(n529), .B(n530), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n458), .B(n381), .ZN(n380) );
  XNOR2_X1 U469 ( .A(n474), .B(n382), .ZN(n381) );
  NAND2_X1 U470 ( .A1(n435), .A2(n356), .ZN(n436) );
  NAND2_X1 U471 ( .A1(n742), .A2(n440), .ZN(n438) );
  XNOR2_X1 U472 ( .A(n656), .B(n401), .ZN(n618) );
  INV_X1 U473 ( .A(KEYINPUT101), .ZN(n401) );
  NAND2_X1 U474 ( .A1(n428), .A2(n583), .ZN(n427) );
  INV_X1 U475 ( .A(KEYINPUT33), .ZN(n394) );
  INV_X1 U476 ( .A(n562), .ZN(n586) );
  AND2_X1 U477 ( .A1(n570), .A2(n375), .ZN(n584) );
  NOR2_X1 U478 ( .A1(n376), .A2(n390), .ZN(n375) );
  INV_X1 U479 ( .A(n574), .ZN(n390) );
  XNOR2_X1 U480 ( .A(n564), .B(KEYINPUT30), .ZN(n376) );
  XNOR2_X1 U481 ( .A(n366), .B(n509), .ZN(n718) );
  XNOR2_X1 U482 ( .A(n508), .B(n449), .ZN(n509) );
  XNOR2_X1 U483 ( .A(n504), .B(n735), .ZN(n366) );
  NOR2_X1 U484 ( .A1(G952), .A2(n743), .ZN(n720) );
  NOR2_X1 U485 ( .A1(n598), .A2(n695), .ZN(n580) );
  XNOR2_X1 U486 ( .A(n374), .B(n362), .ZN(n750) );
  INV_X1 U487 ( .A(KEYINPUT36), .ZN(n389) );
  XNOR2_X1 U488 ( .A(n553), .B(KEYINPUT32), .ZN(n748) );
  XNOR2_X1 U489 ( .A(n600), .B(n599), .ZN(n651) );
  NOR2_X1 U490 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U491 ( .A(n548), .B(KEYINPUT64), .ZN(n406) );
  AND2_X1 U492 ( .A1(n398), .A2(n360), .ZN(n639) );
  XNOR2_X1 U493 ( .A(n404), .B(n403), .ZN(n537) );
  INV_X1 U494 ( .A(KEYINPUT85), .ZN(n403) );
  NAND2_X1 U495 ( .A1(n388), .A2(n358), .ZN(n404) );
  BUF_X1 U496 ( .A(n680), .Z(n405) );
  AND2_X1 U497 ( .A1(n523), .A2(G210), .ZN(n352) );
  XNOR2_X1 U498 ( .A(n492), .B(n491), .ZN(n353) );
  XOR2_X1 U499 ( .A(KEYINPUT95), .B(n498), .Z(n354) );
  XOR2_X1 U500 ( .A(KEYINPUT72), .B(G116), .Z(n355) );
  NOR2_X1 U501 ( .A1(n621), .A2(n434), .ZN(n356) );
  AND2_X1 U502 ( .A1(n386), .A2(n385), .ZN(n357) );
  AND2_X1 U503 ( .A1(n405), .A2(n536), .ZN(n358) );
  OR2_X1 U504 ( .A1(n610), .A2(n609), .ZN(n359) );
  AND2_X1 U505 ( .A1(n570), .A2(n392), .ZN(n360) );
  AND2_X1 U506 ( .A1(n535), .A2(n445), .ZN(n361) );
  INV_X1 U507 ( .A(KEYINPUT104), .ZN(n387) );
  INV_X1 U508 ( .A(KEYINPUT34), .ZN(n432) );
  XOR2_X1 U509 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n362) );
  XNOR2_X1 U510 ( .A(n453), .B(n478), .ZN(n728) );
  XOR2_X1 U511 ( .A(n632), .B(n631), .Z(n363) );
  NAND2_X1 U512 ( .A1(n364), .A2(n378), .ZN(n555) );
  AND2_X1 U513 ( .A1(n365), .A2(n555), .ZN(n559) );
  NOR2_X1 U514 ( .A1(n545), .A2(n544), .ZN(n365) );
  NOR2_X1 U515 ( .A1(n367), .A2(n604), .ZN(n605) );
  XNOR2_X1 U516 ( .A(n603), .B(KEYINPUT76), .ZN(n367) );
  INV_X1 U517 ( .A(n621), .ZN(n369) );
  NAND2_X1 U518 ( .A1(n576), .A2(n575), .ZN(n419) );
  NAND2_X1 U519 ( .A1(n750), .A2(n751), .ZN(n581) );
  NAND2_X1 U520 ( .A1(n617), .A2(n653), .ZN(n374) );
  NOR2_X1 U521 ( .A1(n644), .A2(n748), .ZN(n379) );
  INV_X1 U522 ( .A(n554), .ZN(n377) );
  INV_X1 U523 ( .A(n644), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n379), .A2(n556), .ZN(n557) );
  NAND2_X1 U525 ( .A1(n357), .A2(n383), .ZN(n547) );
  NAND2_X1 U526 ( .A1(n388), .A2(n384), .ZN(n383) );
  INV_X1 U527 ( .A(n550), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n550), .A2(n387), .ZN(n386) );
  INV_X2 U529 ( .A(KEYINPUT68), .ZN(n399) );
  XNOR2_X1 U530 ( .A(n593), .B(n389), .ZN(n594) );
  NAND2_X1 U531 ( .A1(n559), .A2(n558), .ZN(n561) );
  AND2_X1 U532 ( .A1(n605), .A2(n359), .ZN(n391) );
  INV_X1 U533 ( .A(n563), .ZN(n392) );
  XNOR2_X2 U534 ( .A(n393), .B(n353), .ZN(n577) );
  OR2_X2 U535 ( .A1(n707), .A2(G902), .ZN(n393) );
  NAND2_X1 U536 ( .A1(n540), .A2(n589), .ZN(n395) );
  NAND2_X1 U537 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U538 ( .A(n686), .ZN(n397) );
  XNOR2_X2 U539 ( .A(n399), .B(G131), .ZN(n527) );
  XNOR2_X1 U540 ( .A(n591), .B(n463), .ZN(n597) );
  NOR2_X2 U541 ( .A1(n406), .A2(n549), .ZN(n644) );
  XNOR2_X1 U542 ( .A(n581), .B(n410), .ZN(n606) );
  NAND2_X1 U543 ( .A1(n562), .A2(n664), .ZN(n591) );
  XNOR2_X1 U544 ( .A(n499), .B(n521), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n408), .B(n635), .ZN(G60) );
  XNOR2_X1 U546 ( .A(n441), .B(n450), .ZN(n453) );
  XNOR2_X1 U547 ( .A(n409), .B(n706), .ZN(G51) );
  XNOR2_X2 U548 ( .A(n411), .B(n354), .ZN(n676) );
  NAND2_X1 U549 ( .A1(n422), .A2(n412), .ZN(n626) );
  NAND2_X1 U550 ( .A1(n422), .A2(n413), .ZN(n633) );
  NAND2_X1 U551 ( .A1(n422), .A2(n414), .ZN(n704) );
  NAND2_X1 U552 ( .A1(n431), .A2(n361), .ZN(n444) );
  OR2_X1 U553 ( .A1(n431), .A2(n432), .ZN(n428) );
  INV_X1 U554 ( .A(n431), .ZN(n416) );
  NAND2_X1 U555 ( .A1(n417), .A2(n577), .ZN(n578) );
  NOR2_X1 U556 ( .A1(n420), .A2(n651), .ZN(n603) );
  NAND2_X1 U557 ( .A1(n602), .A2(n610), .ZN(n420) );
  AND2_X2 U558 ( .A1(n436), .A2(n423), .ZN(n422) );
  NAND2_X1 U559 ( .A1(n437), .A2(n436), .ZN(n424) );
  INV_X1 U560 ( .A(n622), .ZN(n423) );
  NAND2_X1 U561 ( .A1(n424), .A2(n699), .ZN(n700) );
  NAND2_X1 U562 ( .A1(n426), .A2(n425), .ZN(n446) );
  NAND2_X1 U563 ( .A1(n696), .A2(KEYINPUT34), .ZN(n425) );
  NAND2_X1 U564 ( .A1(n398), .A2(n432), .ZN(n430) );
  OR2_X1 U565 ( .A1(n620), .A2(n440), .ZN(n434) );
  INV_X1 U566 ( .A(n724), .ZN(n435) );
  XNOR2_X2 U567 ( .A(n561), .B(n560), .ZN(n724) );
  AND2_X2 U568 ( .A1(n439), .A2(n438), .ZN(n437) );
  NAND2_X1 U569 ( .A1(n724), .A2(n440), .ZN(n439) );
  INV_X1 U570 ( .A(KEYINPUT2), .ZN(n440) );
  XNOR2_X2 U571 ( .A(n446), .B(KEYINPUT35), .ZN(n546) );
  XNOR2_X1 U572 ( .A(n633), .B(n363), .ZN(n634) );
  XNOR2_X1 U573 ( .A(n702), .B(n448), .ZN(n703) );
  XNOR2_X1 U574 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U575 ( .A(n507), .B(n506), .Z(n449) );
  NAND2_X1 U576 ( .A1(n619), .A2(n662), .ZN(n620) );
  INV_X1 U577 ( .A(KEYINPUT39), .ZN(n571) );
  XNOR2_X1 U578 ( .A(n624), .B(n623), .ZN(n625) );
  INV_X1 U579 ( .A(KEYINPUT78), .ZN(n599) );
  XNOR2_X1 U580 ( .A(n704), .B(n703), .ZN(n705) );
  INV_X1 U581 ( .A(KEYINPUT63), .ZN(n628) );
  XNOR2_X1 U582 ( .A(KEYINPUT60), .B(KEYINPUT120), .ZN(n635) );
  XOR2_X1 U583 ( .A(G128), .B(G143), .Z(n474) );
  XNOR2_X1 U584 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U585 ( .A(n501), .B(n456), .ZN(n458) );
  NAND2_X1 U586 ( .A1(G224), .A2(n743), .ZN(n457) );
  XOR2_X1 U587 ( .A(KEYINPUT74), .B(G107), .Z(n483) );
  XNOR2_X1 U588 ( .A(n459), .B(KEYINPUT77), .ZN(n462) );
  NAND2_X1 U589 ( .A1(n462), .A2(G210), .ZN(n460) );
  NAND2_X1 U590 ( .A1(G214), .A2(n462), .ZN(n664) );
  XOR2_X1 U591 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n463) );
  NAND2_X1 U592 ( .A1(G234), .A2(G237), .ZN(n464) );
  XNOR2_X1 U593 ( .A(n464), .B(KEYINPUT14), .ZN(n466) );
  NAND2_X1 U594 ( .A1(G952), .A2(n466), .ZN(n694) );
  NOR2_X1 U595 ( .A1(n694), .A2(G953), .ZN(n465) );
  XNOR2_X1 U596 ( .A(n465), .B(KEYINPUT89), .ZN(n567) );
  INV_X1 U597 ( .A(n567), .ZN(n469) );
  NAND2_X1 U598 ( .A1(G902), .A2(n466), .ZN(n565) );
  XOR2_X1 U599 ( .A(G898), .B(KEYINPUT90), .Z(n723) );
  NAND2_X1 U600 ( .A1(n723), .A2(G953), .ZN(n467) );
  XOR2_X1 U601 ( .A(KEYINPUT91), .B(n467), .Z(n729) );
  NOR2_X1 U602 ( .A1(n565), .A2(n729), .ZN(n468) );
  NOR2_X1 U603 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U604 ( .A(n470), .B(KEYINPUT92), .ZN(n471) );
  XOR2_X1 U605 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n476) );
  XNOR2_X1 U606 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U607 ( .A(G472), .B(KEYINPUT97), .ZN(n479) );
  XNOR2_X1 U608 ( .A(n563), .B(KEYINPUT103), .ZN(n481) );
  XNOR2_X1 U609 ( .A(n734), .B(G101), .ZN(n490) );
  XNOR2_X1 U610 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U611 ( .A(G104), .B(n485), .Z(n487) );
  NAND2_X1 U612 ( .A1(G227), .A2(n743), .ZN(n486) );
  XNOR2_X1 U613 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U614 ( .A(n488), .B(G140), .Z(n489) );
  XNOR2_X1 U615 ( .A(n490), .B(n489), .ZN(n707) );
  XNOR2_X1 U616 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n492) );
  INV_X1 U617 ( .A(G469), .ZN(n491) );
  NAND2_X1 U618 ( .A1(G234), .A2(n622), .ZN(n494) );
  XNOR2_X1 U619 ( .A(KEYINPUT20), .B(n494), .ZN(n496) );
  NAND2_X1 U620 ( .A1(n496), .A2(G221), .ZN(n495) );
  XNOR2_X1 U621 ( .A(n495), .B(KEYINPUT21), .ZN(n675) );
  NAND2_X1 U622 ( .A1(G217), .A2(n496), .ZN(n497) );
  XNOR2_X1 U623 ( .A(n497), .B(KEYINPUT25), .ZN(n498) );
  XOR2_X1 U624 ( .A(n499), .B(G137), .Z(n500) );
  XNOR2_X1 U625 ( .A(n501), .B(G140), .ZN(n503) );
  XOR2_X1 U626 ( .A(KEYINPUT8), .B(n505), .Z(n512) );
  NAND2_X1 U627 ( .A1(G221), .A2(n512), .ZN(n508) );
  OR2_X1 U628 ( .A1(n675), .A2(n676), .ZN(n679) );
  XOR2_X1 U629 ( .A(KEYINPUT99), .B(G107), .Z(n511) );
  XNOR2_X1 U630 ( .A(G116), .B(G122), .ZN(n510) );
  XNOR2_X1 U631 ( .A(n511), .B(n510), .ZN(n516) );
  XOR2_X1 U632 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n514) );
  NAND2_X1 U633 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U634 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U635 ( .A(n516), .B(n515), .ZN(n518) );
  XNOR2_X1 U636 ( .A(n517), .B(n518), .ZN(n715) );
  NOR2_X1 U637 ( .A1(G902), .A2(n715), .ZN(n520) );
  XNOR2_X1 U638 ( .A(KEYINPUT100), .B(G478), .ZN(n519) );
  XNOR2_X1 U639 ( .A(n520), .B(n519), .ZN(n538) );
  XNOR2_X1 U640 ( .A(n521), .B(n522), .ZN(n530) );
  NAND2_X1 U641 ( .A1(G214), .A2(n523), .ZN(n524) );
  XNOR2_X1 U642 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U643 ( .A(n526), .B(KEYINPUT98), .Z(n529) );
  XNOR2_X1 U644 ( .A(n527), .B(n735), .ZN(n528) );
  NOR2_X1 U645 ( .A1(G902), .A2(n630), .ZN(n532) );
  XNOR2_X1 U646 ( .A(KEYINPUT13), .B(G475), .ZN(n531) );
  XNOR2_X1 U647 ( .A(n532), .B(n531), .ZN(n539) );
  INV_X1 U648 ( .A(n539), .ZN(n534) );
  NOR2_X1 U649 ( .A1(n538), .A2(n534), .ZN(n583) );
  NOR2_X1 U650 ( .A1(KEYINPUT86), .A2(n533), .ZN(n545) );
  NAND2_X1 U651 ( .A1(n538), .A2(n534), .ZN(n667) );
  INV_X1 U652 ( .A(n667), .ZN(n535) );
  INV_X1 U653 ( .A(n405), .ZN(n614) );
  INV_X1 U654 ( .A(n589), .ZN(n536) );
  NOR2_X1 U655 ( .A1(n676), .A2(n537), .ZN(n636) );
  NAND2_X1 U656 ( .A1(n539), .A2(n538), .ZN(n650) );
  INV_X1 U657 ( .A(n650), .ZN(n653) );
  NOR2_X1 U658 ( .A1(n653), .A2(n618), .ZN(n669) );
  INV_X1 U659 ( .A(n669), .ZN(n607) );
  NAND2_X1 U660 ( .A1(n563), .A2(n540), .ZN(n686) );
  NOR2_X1 U661 ( .A1(n657), .A2(n639), .ZN(n541) );
  NOR2_X1 U662 ( .A1(n601), .A2(n541), .ZN(n542) );
  INV_X1 U663 ( .A(n676), .ZN(n549) );
  NAND2_X1 U664 ( .A1(n547), .A2(n392), .ZN(n548) );
  NOR2_X1 U665 ( .A1(n589), .A2(n550), .ZN(n551) );
  NAND2_X1 U666 ( .A1(n676), .A2(n551), .ZN(n552) );
  NOR2_X1 U667 ( .A1(n552), .A2(n405), .ZN(n553) );
  NAND2_X1 U668 ( .A1(n546), .A2(KEYINPUT86), .ZN(n556) );
  NAND2_X1 U669 ( .A1(n557), .A2(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U670 ( .A1(n664), .A2(n563), .ZN(n564) );
  NOR2_X1 U671 ( .A1(G900), .A2(n565), .ZN(n566) );
  NAND2_X1 U672 ( .A1(n566), .A2(G953), .ZN(n568) );
  NAND2_X1 U673 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U674 ( .A(n569), .B(KEYINPUT80), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n676), .A2(n574), .ZN(n587) );
  INV_X1 U676 ( .A(n587), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n578), .B(KEYINPUT106), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n665), .A2(n664), .ZN(n668) );
  XNOR2_X1 U679 ( .A(n579), .B(KEYINPUT41), .ZN(n695) );
  XOR2_X1 U680 ( .A(KEYINPUT42), .B(n580), .Z(n751) );
  NAND2_X1 U681 ( .A1(KEYINPUT47), .A2(n669), .ZN(n582) );
  NAND2_X1 U682 ( .A1(n582), .A2(KEYINPUT81), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U684 ( .A1(n586), .A2(n585), .ZN(n649) );
  NOR2_X1 U685 ( .A1(n650), .A2(n587), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U687 ( .A(n612), .ZN(n592) );
  NOR2_X1 U688 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U689 ( .A1(n405), .A2(n594), .ZN(n660) );
  NOR2_X1 U690 ( .A1(n649), .A2(n660), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n596), .A2(n595), .ZN(n604) );
  INV_X1 U692 ( .A(KEYINPUT47), .ZN(n610) );
  NOR2_X1 U693 ( .A1(KEYINPUT81), .A2(n607), .ZN(n608) );
  NOR2_X1 U694 ( .A1(n651), .A2(n608), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n612), .A2(n664), .ZN(n613) );
  NOR2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(KEYINPUT43), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n562), .A2(n616), .ZN(n663) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n662) );
  XOR2_X1 U700 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n623) );
  XNOR2_X1 U701 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(G57) );
  XNOR2_X1 U703 ( .A(KEYINPUT119), .B(KEYINPUT65), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT59), .ZN(n631) );
  XOR2_X1 U705 ( .A(G101), .B(n636), .Z(G3) );
  NAND2_X1 U706 ( .A1(n639), .A2(n653), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT108), .ZN(n638) );
  XNOR2_X1 U708 ( .A(G104), .B(n638), .ZN(G6) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U710 ( .A1(n639), .A2(n656), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U712 ( .A(G107), .B(KEYINPUT109), .Z(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G9) );
  XOR2_X1 U714 ( .A(n644), .B(G110), .Z(n645) );
  XNOR2_X1 U715 ( .A(KEYINPUT110), .B(n645), .ZN(G12) );
  XOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .Z(n648) );
  INV_X1 U717 ( .A(n651), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n656), .A2(n646), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(G30) );
  XOR2_X1 U720 ( .A(G143), .B(n649), .Z(G45) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U722 ( .A(G146), .B(n652), .Z(G48) );
  XOR2_X1 U723 ( .A(G113), .B(KEYINPUT111), .Z(n655) );
  NAND2_X1 U724 ( .A1(n657), .A2(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n658), .B(KEYINPUT112), .ZN(n659) );
  XNOR2_X1 U728 ( .A(G116), .B(n659), .ZN(G18) );
  XNOR2_X1 U729 ( .A(G125), .B(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U731 ( .A(G134), .B(n662), .ZN(G36) );
  XOR2_X1 U732 ( .A(G140), .B(n663), .Z(G42) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT115), .B(n670), .Z(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n673), .B(KEYINPUT116), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n400), .A2(n674), .ZN(n691) );
  XOR2_X1 U740 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n678) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n678), .B(n677), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n405), .A2(n679), .ZN(n681) );
  XOR2_X1 U744 ( .A(KEYINPUT50), .B(n681), .Z(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U746 ( .A1(n684), .A2(n392), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT114), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(KEYINPUT51), .B(n688), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n695), .A2(n689), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n692), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U754 ( .A1(n400), .A2(n695), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U756 ( .A1(n700), .A2(G953), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n701), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U758 ( .A(KEYINPUT56), .B(KEYINPUT117), .Z(n706) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n709) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT118), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(n712) );
  NAND2_X1 U762 ( .A1(n710), .A2(G469), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n720), .A2(n713), .ZN(G54) );
  NAND2_X1 U765 ( .A1(G478), .A2(n710), .ZN(n714) );
  NAND2_X1 U766 ( .A1(G217), .A2(n710), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U768 ( .A1(n720), .A2(n719), .ZN(G66) );
  NAND2_X1 U769 ( .A1(G953), .A2(G224), .ZN(n721) );
  XOR2_X1 U770 ( .A(KEYINPUT61), .B(n721), .Z(n722) );
  NOR2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U772 ( .A1(G953), .A2(n724), .ZN(n725) );
  XOR2_X1 U773 ( .A(KEYINPUT121), .B(n725), .Z(n726) );
  NOR2_X1 U774 ( .A1(n727), .A2(n726), .ZN(n733) );
  XNOR2_X1 U775 ( .A(n728), .B(G107), .ZN(n730) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U777 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  XNOR2_X1 U778 ( .A(n733), .B(n732), .ZN(G69) );
  XOR2_X1 U779 ( .A(n734), .B(n735), .Z(n736) );
  XNOR2_X1 U780 ( .A(KEYINPUT123), .B(n736), .ZN(n741) );
  XNOR2_X1 U781 ( .A(G227), .B(n741), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n737), .A2(G900), .ZN(n738) );
  XOR2_X1 U783 ( .A(KEYINPUT124), .B(n738), .Z(n739) );
  NOR2_X1 U784 ( .A1(n743), .A2(n739), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(KEYINPUT125), .ZN(n746) );
  XNOR2_X1 U786 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U787 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U788 ( .A1(n746), .A2(n745), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G122), .B(KEYINPUT126), .ZN(n747) );
  XOR2_X1 U790 ( .A(n747), .B(n546), .Z(G24) );
  XNOR2_X1 U791 ( .A(G119), .B(KEYINPUT127), .ZN(n749) );
  XNOR2_X1 U792 ( .A(n749), .B(n748), .ZN(G21) );
  XNOR2_X1 U793 ( .A(G131), .B(n750), .ZN(G33) );
  XNOR2_X1 U794 ( .A(n751), .B(G137), .ZN(G39) );
endmodule

