

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780;

  XNOR2_X1 U382 ( .A(G116), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X2 U383 ( .A(n770), .B(n439), .ZN(n446) );
  XNOR2_X2 U384 ( .A(n434), .B(n361), .ZN(n525) );
  BUF_X4 U385 ( .A(n544), .Z(n400) );
  NOR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n518) );
  AND2_X1 U387 ( .A1(n411), .A2(n630), .ZN(n631) );
  NOR2_X1 U388 ( .A1(n561), .A2(n562), .ZN(n700) );
  XNOR2_X2 U389 ( .A(n530), .B(n529), .ZN(n597) );
  XNOR2_X2 U390 ( .A(n655), .B(n505), .ZN(n680) );
  OR2_X2 U391 ( .A1(n664), .A2(n427), .ZN(n416) );
  AND2_X2 U392 ( .A1(n664), .A2(n448), .ZN(n399) );
  XNOR2_X2 U393 ( .A(n446), .B(n445), .ZN(n664) );
  XNOR2_X2 U394 ( .A(n525), .B(n363), .ZN(n770) );
  NOR2_X1 U395 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U396 ( .A1(n700), .A2(n696), .ZN(n565) );
  XNOR2_X2 U397 ( .A(n585), .B(KEYINPUT1), .ZN(n544) );
  NAND2_X1 U398 ( .A1(n637), .A2(n419), .ZN(n418) );
  NAND2_X1 U399 ( .A1(n430), .A2(n420), .ZN(n419) );
  AND2_X1 U400 ( .A1(n537), .A2(n539), .ZN(n695) );
  NOR2_X1 U401 ( .A1(n625), .A2(n704), .ZN(n617) );
  NOR2_X1 U402 ( .A1(n597), .A2(n557), .ZN(n734) );
  AND2_X1 U403 ( .A1(n394), .A2(n392), .ZN(n391) );
  NAND2_X1 U404 ( .A1(n385), .A2(n383), .ZN(n592) );
  XNOR2_X1 U405 ( .A(n602), .B(n612), .ZN(n739) );
  AND2_X1 U406 ( .A1(n416), .A2(n405), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n435), .B(G953), .ZN(n500) );
  XNOR2_X1 U408 ( .A(n415), .B(G119), .ZN(n434) );
  XNOR2_X1 U409 ( .A(n664), .B(n666), .ZN(n667) );
  XNOR2_X2 U410 ( .A(n485), .B(n484), .ZN(n498) );
  XNOR2_X2 U411 ( .A(n460), .B(KEYINPUT0), .ZN(n548) );
  INV_X1 U412 ( .A(n382), .ZN(n381) );
  XOR2_X1 U413 ( .A(KEYINPUT75), .B(G137), .Z(n496) );
  XNOR2_X1 U414 ( .A(KEYINPUT72), .B(G101), .ZN(n522) );
  AND2_X1 U415 ( .A1(n403), .A2(n371), .ZN(n402) );
  NAND2_X1 U416 ( .A1(n423), .A2(KEYINPUT68), .ZN(n403) );
  NAND2_X1 U417 ( .A1(n543), .A2(KEYINPUT68), .ZN(n404) );
  NAND2_X1 U418 ( .A1(n402), .A2(n542), .ZN(n376) );
  NAND2_X1 U419 ( .A1(n404), .A2(KEYINPUT93), .ZN(n375) );
  NAND2_X1 U420 ( .A1(n380), .A2(n379), .ZN(n378) );
  NAND2_X1 U421 ( .A1(n404), .A2(n542), .ZN(n379) );
  NAND2_X1 U422 ( .A1(n402), .A2(KEYINPUT93), .ZN(n380) );
  NAND2_X1 U423 ( .A1(n541), .A2(n540), .ZN(n382) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n464) );
  XNOR2_X1 U425 ( .A(n398), .B(n369), .ZN(n622) );
  NAND2_X1 U426 ( .A1(n393), .A2(KEYINPUT108), .ZN(n392) );
  INV_X1 U427 ( .A(n723), .ZN(n393) );
  INV_X1 U428 ( .A(n591), .ZN(n546) );
  XOR2_X1 U429 ( .A(G131), .B(G140), .Z(n499) );
  INV_X1 U430 ( .A(G128), .ZN(n437) );
  NAND2_X1 U431 ( .A1(n633), .A2(n428), .ZN(n427) );
  INV_X1 U432 ( .A(n448), .ZN(n428) );
  NOR2_X1 U433 ( .A1(n582), .A2(n362), .ZN(n583) );
  NOR2_X2 U434 ( .A1(n725), .A2(n726), .ZN(n723) );
  XNOR2_X1 U435 ( .A(n526), .B(n527), .ZN(n397) );
  XOR2_X1 U436 ( .A(KEYINPUT74), .B(KEYINPUT8), .Z(n480) );
  XNOR2_X1 U437 ( .A(G128), .B(G140), .ZN(n508) );
  XNOR2_X1 U438 ( .A(n407), .B(KEYINPUT24), .ZN(n509) );
  INV_X1 U439 ( .A(KEYINPUT23), .ZN(n407) );
  XNOR2_X1 U440 ( .A(G119), .B(G137), .ZN(n507) );
  XOR2_X1 U441 ( .A(KEYINPUT10), .B(n462), .Z(n654) );
  XNOR2_X1 U442 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X1 U443 ( .A(KEYINPUT82), .B(KEYINPUT17), .ZN(n442) );
  NOR2_X1 U444 ( .A1(n613), .A2(n739), .ZN(n616) );
  BUF_X1 U445 ( .A(n500), .Z(n656) );
  NAND2_X1 U446 ( .A1(n382), .A2(n374), .ZN(n373) );
  NAND2_X1 U447 ( .A1(n381), .A2(n378), .ZN(n377) );
  NAND2_X1 U448 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U449 ( .A1(n778), .A2(n422), .ZN(n424) );
  AND2_X1 U450 ( .A1(n553), .A2(KEYINPUT68), .ZN(n422) );
  XOR2_X1 U451 ( .A(G146), .B(G131), .Z(n520) );
  XNOR2_X1 U452 ( .A(G113), .B(G104), .ZN(n465) );
  XNOR2_X1 U453 ( .A(G143), .B(G122), .ZN(n463) );
  AND2_X1 U454 ( .A1(n431), .A2(n421), .ZN(n420) );
  INV_X1 U455 ( .A(KEYINPUT89), .ZN(n421) );
  NAND2_X1 U456 ( .A1(n634), .A2(KEYINPUT2), .ZN(n431) );
  XNOR2_X1 U457 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U458 ( .A1(G234), .A2(G237), .ZN(n452) );
  XOR2_X1 U459 ( .A(KEYINPUT14), .B(KEYINPUT97), .Z(n453) );
  INV_X1 U460 ( .A(G237), .ZN(n447) );
  NOR2_X1 U461 ( .A1(n739), .A2(n738), .ZN(n744) );
  XNOR2_X1 U462 ( .A(n547), .B(KEYINPUT33), .ZN(n737) );
  NAND2_X1 U463 ( .A1(n391), .A2(n389), .ZN(n547) );
  AND2_X1 U464 ( .A1(n546), .A2(n390), .ZN(n389) );
  NAND2_X1 U465 ( .A1(n634), .A2(n448), .ZN(n429) );
  NAND2_X1 U466 ( .A1(n364), .A2(n414), .ZN(n590) );
  INV_X1 U467 ( .A(n725), .ZN(n414) );
  XNOR2_X1 U468 ( .A(G122), .B(KEYINPUT9), .ZN(n476) );
  XOR2_X1 U469 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n477) );
  INV_X1 U470 ( .A(G134), .ZN(n484) );
  BUF_X1 U471 ( .A(n737), .Z(n755) );
  XNOR2_X1 U472 ( .A(n412), .B(KEYINPUT109), .ZN(n627) );
  NAND2_X1 U473 ( .A1(n413), .A2(n700), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n591), .A2(n590), .ZN(n413) );
  NOR2_X1 U475 ( .A1(n600), .A2(n396), .ZN(n395) );
  INV_X1 U476 ( .A(n601), .ZN(n396) );
  XNOR2_X1 U477 ( .A(n592), .B(KEYINPUT19), .ZN(n588) );
  XNOR2_X1 U478 ( .A(n647), .B(n646), .ZN(n648) );
  AND2_X1 U479 ( .A1(n512), .A2(G221), .ZN(n408) );
  XOR2_X1 U480 ( .A(G146), .B(KEYINPUT99), .Z(n502) );
  NOR2_X1 U481 ( .A1(n656), .A2(G952), .ZN(n683) );
  XNOR2_X1 U482 ( .A(n621), .B(KEYINPUT42), .ZN(n779) );
  AND2_X1 U483 ( .A1(n588), .A2(n620), .ZN(n701) );
  INV_X1 U484 ( .A(n700), .ZN(n704) );
  AND2_X1 U485 ( .A1(n416), .A2(n429), .ZN(n360) );
  XOR2_X1 U486 ( .A(G113), .B(KEYINPUT76), .Z(n361) );
  AND2_X1 U487 ( .A1(n581), .A2(n580), .ZN(n362) );
  NAND2_X1 U488 ( .A1(n360), .A2(n387), .ZN(n602) );
  XOR2_X1 U489 ( .A(KEYINPUT16), .B(G122), .Z(n363) );
  AND2_X1 U490 ( .A1(n726), .A2(n601), .ZN(n364) );
  AND2_X1 U491 ( .A1(n631), .A2(n634), .ZN(n365) );
  XOR2_X1 U492 ( .A(n599), .B(n598), .Z(n366) );
  AND2_X1 U493 ( .A1(n608), .A2(KEYINPUT47), .ZN(n367) );
  AND2_X1 U494 ( .A1(n723), .A2(n545), .ZN(n368) );
  NAND2_X1 U495 ( .A1(n429), .A2(n426), .ZN(n425) );
  INV_X1 U496 ( .A(KEYINPUT94), .ZN(n405) );
  INV_X1 U497 ( .A(n543), .ZN(n423) );
  XOR2_X1 U498 ( .A(KEYINPUT65), .B(KEYINPUT46), .Z(n369) );
  XOR2_X1 U499 ( .A(n639), .B(n638), .Z(n370) );
  NAND2_X1 U500 ( .A1(n554), .A2(KEYINPUT44), .ZN(n371) );
  NAND2_X1 U501 ( .A1(n377), .A2(n373), .ZN(n401) );
  AND2_X1 U502 ( .A1(n710), .A2(n432), .ZN(n610) );
  XNOR2_X2 U503 ( .A(n372), .B(KEYINPUT45), .ZN(n713) );
  NAND2_X1 U504 ( .A1(n576), .A2(n577), .ZN(n372) );
  NAND2_X1 U505 ( .A1(n406), .A2(n384), .ZN(n383) );
  NAND2_X1 U506 ( .A1(n386), .A2(KEYINPUT94), .ZN(n385) );
  NAND2_X1 U507 ( .A1(n406), .A2(n416), .ZN(n386) );
  INV_X1 U508 ( .A(n399), .ZN(n387) );
  XNOR2_X1 U509 ( .A(n388), .B(n397), .ZN(n647) );
  XNOR2_X2 U510 ( .A(n388), .B(n499), .ZN(n655) );
  XNOR2_X2 U511 ( .A(n498), .B(n497), .ZN(n388) );
  NAND2_X1 U512 ( .A1(n400), .A2(n723), .ZN(n557) );
  NAND2_X1 U513 ( .A1(n544), .A2(n368), .ZN(n390) );
  OR2_X2 U514 ( .A1(n544), .A2(n545), .ZN(n394) );
  NAND2_X1 U515 ( .A1(n366), .A2(n395), .ZN(n613) );
  NAND2_X1 U516 ( .A1(n780), .A2(n779), .ZN(n398) );
  NAND2_X1 U517 ( .A1(n707), .A2(n689), .ZN(n567) );
  XNOR2_X2 U518 ( .A(n560), .B(n559), .ZN(n707) );
  XNOR2_X1 U519 ( .A(n536), .B(n535), .ZN(n663) );
  XNOR2_X1 U520 ( .A(n494), .B(KEYINPUT22), .ZN(n537) );
  NOR2_X1 U521 ( .A1(n399), .A2(n425), .ZN(n406) );
  NAND2_X1 U522 ( .A1(n537), .A2(n534), .ZN(n536) );
  NAND2_X1 U523 ( .A1(n401), .A2(n424), .ZN(n577) );
  NOR2_X1 U524 ( .A1(n671), .A2(G902), .ZN(n517) );
  XNOR2_X1 U525 ( .A(n409), .B(n408), .ZN(n671) );
  XNOR2_X1 U526 ( .A(n654), .B(n410), .ZN(n409) );
  XNOR2_X1 U527 ( .A(n510), .B(n511), .ZN(n410) );
  INV_X1 U528 ( .A(n631), .ZN(n716) );
  XNOR2_X1 U529 ( .A(n624), .B(KEYINPUT48), .ZN(n411) );
  AND2_X2 U530 ( .A1(n713), .A2(n631), .ZN(n720) );
  XNOR2_X2 U531 ( .A(n417), .B(n437), .ZN(n485) );
  XNOR2_X2 U532 ( .A(G143), .B(KEYINPUT66), .ZN(n417) );
  XNOR2_X2 U533 ( .A(n418), .B(KEYINPUT67), .ZN(n674) );
  XNOR2_X2 U534 ( .A(n552), .B(KEYINPUT35), .ZN(n778) );
  INV_X1 U535 ( .A(n738), .ZN(n426) );
  NAND2_X1 U536 ( .A1(n713), .A2(n365), .ZN(n430) );
  NOR2_X1 U537 ( .A1(n609), .A2(n367), .ZN(n432) );
  XOR2_X1 U538 ( .A(n643), .B(KEYINPUT71), .Z(n433) );
  INV_X1 U539 ( .A(KEYINPUT5), .ZN(n521) );
  INV_X1 U540 ( .A(KEYINPUT108), .ZN(n545) );
  XNOR2_X1 U541 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U542 ( .A(KEYINPUT30), .ZN(n598) );
  XNOR2_X1 U543 ( .A(n524), .B(n523), .ZN(n527) );
  BUF_X1 U544 ( .A(n713), .Z(n714) );
  XNOR2_X1 U545 ( .A(KEYINPUT13), .B(G475), .ZN(n473) );
  XNOR2_X1 U546 ( .A(n474), .B(n473), .ZN(n563) );
  INV_X1 U547 ( .A(n683), .ZN(n641) );
  INV_X1 U548 ( .A(KEYINPUT63), .ZN(n651) );
  INV_X1 U549 ( .A(KEYINPUT64), .ZN(n435) );
  NAND2_X1 U550 ( .A1(n500), .A2(G224), .ZN(n436) );
  XNOR2_X1 U551 ( .A(KEYINPUT73), .B(KEYINPUT4), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n436), .B(n495), .ZN(n438) );
  XNOR2_X1 U553 ( .A(n485), .B(n438), .ZN(n439) );
  XNOR2_X1 U554 ( .A(G107), .B(G104), .ZN(n441) );
  XNOR2_X1 U555 ( .A(KEYINPUT80), .B(G110), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n441), .B(n440), .ZN(n772) );
  XNOR2_X1 U557 ( .A(n772), .B(n522), .ZN(n504) );
  XNOR2_X1 U558 ( .A(n442), .B(KEYINPUT18), .ZN(n443) );
  XNOR2_X1 U559 ( .A(n461), .B(n443), .ZN(n444) );
  XNOR2_X1 U560 ( .A(n504), .B(n444), .ZN(n445) );
  XNOR2_X1 U561 ( .A(KEYINPUT15), .B(G902), .ZN(n633) );
  INV_X1 U562 ( .A(n633), .ZN(n634) );
  INV_X1 U563 ( .A(G902), .ZN(n528) );
  NAND2_X1 U564 ( .A1(n528), .A2(n447), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n449), .A2(G210), .ZN(n448) );
  NAND2_X1 U566 ( .A1(n449), .A2(G214), .ZN(n451) );
  INV_X1 U567 ( .A(KEYINPUT96), .ZN(n450) );
  XNOR2_X1 U568 ( .A(n451), .B(n450), .ZN(n738) );
  NAND2_X1 U569 ( .A1(G952), .A2(n454), .ZN(n752) );
  NOR2_X1 U570 ( .A1(n752), .A2(G953), .ZN(n582) );
  INV_X1 U571 ( .A(n582), .ZN(n458) );
  NAND2_X1 U572 ( .A1(n454), .A2(G902), .ZN(n455) );
  XOR2_X1 U573 ( .A(KEYINPUT98), .B(n455), .Z(n581) );
  INV_X1 U574 ( .A(G898), .ZN(n456) );
  AND2_X1 U575 ( .A1(n456), .A2(G953), .ZN(n774) );
  NAND2_X1 U576 ( .A1(n581), .A2(n774), .ZN(n457) );
  NAND2_X1 U577 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U578 ( .A1(n588), .A2(n459), .ZN(n460) );
  INV_X1 U579 ( .A(n461), .ZN(n462) );
  XOR2_X1 U580 ( .A(n654), .B(n499), .Z(n472) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U582 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U583 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n468) );
  NAND2_X1 U584 ( .A1(G214), .A2(n518), .ZN(n467) );
  XNOR2_X1 U585 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U586 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U587 ( .A(n472), .B(n471), .ZN(n639) );
  NOR2_X1 U588 ( .A1(G902), .A2(n639), .ZN(n474) );
  INV_X1 U589 ( .A(n563), .ZN(n562) );
  XNOR2_X1 U590 ( .A(G116), .B(G107), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n475), .B(KEYINPUT7), .ZN(n479) );
  XNOR2_X1 U592 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U593 ( .A(n479), .B(n478), .Z(n483) );
  NAND2_X1 U594 ( .A1(n500), .A2(G234), .ZN(n481) );
  XNOR2_X1 U595 ( .A(n481), .B(n480), .ZN(n512) );
  NAND2_X1 U596 ( .A1(G217), .A2(n512), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n483), .B(n482), .ZN(n487) );
  INV_X1 U598 ( .A(n498), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n487), .B(n486), .ZN(n675) );
  NOR2_X1 U600 ( .A1(G902), .A2(n675), .ZN(n488) );
  XNOR2_X1 U601 ( .A(G478), .B(n488), .ZN(n564) );
  NAND2_X1 U602 ( .A1(n562), .A2(n564), .ZN(n618) );
  NAND2_X1 U603 ( .A1(n633), .A2(G234), .ZN(n489) );
  XNOR2_X1 U604 ( .A(n489), .B(KEYINPUT20), .ZN(n513) );
  NAND2_X1 U605 ( .A1(n513), .A2(G221), .ZN(n490) );
  XNOR2_X1 U606 ( .A(KEYINPUT21), .B(n490), .ZN(n725) );
  NOR2_X1 U607 ( .A1(n618), .A2(n725), .ZN(n492) );
  INV_X1 U608 ( .A(KEYINPUT106), .ZN(n491) );
  XNOR2_X1 U609 ( .A(n492), .B(n491), .ZN(n493) );
  NOR2_X2 U610 ( .A1(n548), .A2(n493), .ZN(n494) );
  XNOR2_X1 U611 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U612 ( .A1(n656), .A2(G227), .ZN(n501) );
  XNOR2_X1 U613 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U614 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U615 ( .A1(n680), .A2(n528), .ZN(n506) );
  XNOR2_X2 U616 ( .A(n506), .B(G469), .ZN(n585) );
  XNOR2_X1 U617 ( .A(n507), .B(G110), .ZN(n511) );
  XNOR2_X1 U618 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U619 ( .A1(n513), .A2(G217), .ZN(n515) );
  XNOR2_X1 U620 ( .A(KEYINPUT25), .B(KEYINPUT81), .ZN(n514) );
  XNOR2_X1 U621 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X2 U622 ( .A(n517), .B(n516), .ZN(n726) );
  NAND2_X1 U623 ( .A1(n400), .A2(n726), .ZN(n533) );
  NAND2_X1 U624 ( .A1(n518), .A2(G210), .ZN(n519) );
  XNOR2_X1 U625 ( .A(n520), .B(n519), .ZN(n524) );
  INV_X1 U626 ( .A(n525), .ZN(n526) );
  NAND2_X1 U627 ( .A1(n647), .A2(n528), .ZN(n530) );
  INV_X1 U628 ( .A(G472), .ZN(n529) );
  INV_X1 U629 ( .A(KEYINPUT6), .ZN(n531) );
  XNOR2_X1 U630 ( .A(n597), .B(n531), .ZN(n591) );
  XNOR2_X1 U631 ( .A(n591), .B(KEYINPUT83), .ZN(n532) );
  NOR2_X1 U632 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U633 ( .A(KEYINPUT69), .B(KEYINPUT32), .ZN(n535) );
  INV_X1 U634 ( .A(n663), .ZN(n541) );
  NAND2_X1 U635 ( .A1(n726), .A2(n597), .ZN(n538) );
  NOR2_X1 U636 ( .A1(n400), .A2(n538), .ZN(n539) );
  INV_X1 U637 ( .A(n695), .ZN(n540) );
  INV_X1 U638 ( .A(KEYINPUT93), .ZN(n542) );
  INV_X1 U639 ( .A(KEYINPUT44), .ZN(n553) );
  NAND2_X1 U640 ( .A1(n553), .A2(KEYINPUT92), .ZN(n543) );
  INV_X1 U641 ( .A(n548), .ZN(n558) );
  NAND2_X1 U642 ( .A1(n737), .A2(n558), .ZN(n550) );
  INV_X1 U643 ( .A(KEYINPUT34), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n550), .B(n549), .ZN(n551) );
  NOR2_X1 U645 ( .A1(n562), .A2(n564), .ZN(n604) );
  NAND2_X1 U646 ( .A1(n551), .A2(n604), .ZN(n552) );
  INV_X1 U647 ( .A(KEYINPUT68), .ZN(n554) );
  NAND2_X1 U648 ( .A1(n778), .A2(KEYINPUT44), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n585), .A2(n723), .ZN(n600) );
  INV_X1 U650 ( .A(n597), .ZN(n555) );
  NOR2_X1 U651 ( .A1(n600), .A2(n555), .ZN(n556) );
  NAND2_X1 U652 ( .A1(n558), .A2(n556), .ZN(n689) );
  NAND2_X1 U653 ( .A1(n558), .A2(n734), .ZN(n560) );
  XOR2_X1 U654 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n559) );
  INV_X1 U655 ( .A(n564), .ZN(n561) );
  NOR2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n696) );
  XNOR2_X1 U657 ( .A(KEYINPUT105), .B(n565), .ZN(n743) );
  INV_X1 U658 ( .A(n743), .ZN(n596) );
  XOR2_X1 U659 ( .A(KEYINPUT87), .B(n596), .Z(n578) );
  INV_X1 U660 ( .A(n578), .ZN(n566) );
  NAND2_X1 U661 ( .A1(n567), .A2(n566), .ZN(n571) );
  NOR2_X1 U662 ( .A1(n400), .A2(n726), .ZN(n568) );
  AND2_X1 U663 ( .A1(n568), .A2(n591), .ZN(n569) );
  NAND2_X1 U664 ( .A1(n537), .A2(n569), .ZN(n685) );
  NAND2_X1 U665 ( .A1(n571), .A2(n685), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n572), .B(KEYINPUT107), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n573), .A2(n574), .ZN(n575) );
  XNOR2_X1 U668 ( .A(n575), .B(KEYINPUT91), .ZN(n576) );
  NOR2_X1 U669 ( .A1(KEYINPUT47), .A2(n578), .ZN(n579) );
  XNOR2_X1 U670 ( .A(KEYINPUT78), .B(n579), .ZN(n589) );
  NOR2_X1 U671 ( .A1(n656), .A2(G900), .ZN(n580) );
  XOR2_X1 U672 ( .A(KEYINPUT84), .B(n583), .Z(n601) );
  NOR2_X1 U673 ( .A1(n597), .A2(n590), .ZN(n584) );
  XOR2_X1 U674 ( .A(KEYINPUT28), .B(n584), .Z(n587) );
  INV_X1 U675 ( .A(n585), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n587), .A2(n586), .ZN(n620) );
  NAND2_X1 U677 ( .A1(n589), .A2(n701), .ZN(n611) );
  INV_X1 U678 ( .A(n592), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n627), .A2(n593), .ZN(n594) );
  XOR2_X1 U680 ( .A(n594), .B(KEYINPUT36), .Z(n595) );
  NAND2_X1 U681 ( .A1(n595), .A2(n400), .ZN(n710) );
  NAND2_X1 U682 ( .A1(n596), .A2(KEYINPUT47), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n597), .A2(n738), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n613), .A2(n602), .ZN(n603) );
  XNOR2_X1 U685 ( .A(n603), .B(KEYINPUT110), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n699) );
  NAND2_X1 U687 ( .A1(n606), .A2(n699), .ZN(n607) );
  XNOR2_X1 U688 ( .A(KEYINPUT86), .B(n607), .ZN(n609) );
  INV_X1 U689 ( .A(n701), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n623) );
  XNOR2_X1 U691 ( .A(KEYINPUT38), .B(KEYINPUT79), .ZN(n612) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(KEYINPUT90), .Z(n614) );
  XNOR2_X1 U693 ( .A(KEYINPUT39), .B(n614), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n616), .B(n615), .ZN(n625) );
  XOR2_X1 U695 ( .A(KEYINPUT40), .B(n617), .Z(n780) );
  INV_X1 U696 ( .A(n618), .ZN(n741) );
  NAND2_X1 U697 ( .A1(n744), .A2(n741), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT41), .ZN(n754) );
  NAND2_X1 U699 ( .A1(n620), .A2(n754), .ZN(n621) );
  INV_X1 U700 ( .A(n696), .ZN(n706) );
  NOR2_X1 U701 ( .A1(n625), .A2(n706), .ZN(n711) );
  NOR2_X1 U702 ( .A1(n738), .A2(n400), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  AND2_X1 U705 ( .A1(n629), .A2(n602), .ZN(n653) );
  NOR2_X1 U706 ( .A1(n711), .A2(n653), .ZN(n630) );
  INV_X1 U707 ( .A(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n634), .A2(KEYINPUT89), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n635), .A2(n632), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n720), .A2(n636), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n674), .A2(G475), .ZN(n640) );
  XOR2_X1 U712 ( .A(KEYINPUT70), .B(KEYINPUT59), .Z(n638) );
  XNOR2_X1 U713 ( .A(n640), .B(n370), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U715 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n644), .B(n433), .ZN(G60) );
  NAND2_X1 U717 ( .A1(n674), .A2(G472), .ZN(n649) );
  XOR2_X1 U718 ( .A(KEYINPUT95), .B(KEYINPUT111), .Z(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(KEYINPUT62), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X2 U721 ( .A1(n650), .A2(n683), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(G57) );
  XOR2_X1 U723 ( .A(n653), .B(G140), .Z(G42) );
  XOR2_X1 U724 ( .A(n655), .B(n654), .Z(n658) );
  XNOR2_X1 U725 ( .A(n716), .B(n658), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n662) );
  XNOR2_X1 U727 ( .A(G227), .B(n658), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n659), .A2(G900), .ZN(n660) );
  NAND2_X1 U729 ( .A1(G953), .A2(n660), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(G72) );
  XOR2_X1 U731 ( .A(n663), .B(G119), .Z(G21) );
  NAND2_X1 U732 ( .A1(n674), .A2(G210), .ZN(n668) );
  XNOR2_X1 U733 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n665) );
  XOR2_X1 U734 ( .A(n665), .B(KEYINPUT55), .Z(n666) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U736 ( .A1(n669), .A2(n683), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U738 ( .A(n674), .Z(n678) );
  NAND2_X1 U739 ( .A1(n678), .A2(G217), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n671), .B(n672), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n673), .A2(n683), .ZN(G66) );
  NAND2_X1 U742 ( .A1(n678), .A2(G478), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n677), .A2(n683), .ZN(G63) );
  NAND2_X1 U745 ( .A1(n678), .A2(G469), .ZN(n682) );
  XNOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n682), .B(n681), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(G54) );
  XNOR2_X1 U750 ( .A(G101), .B(KEYINPUT112), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(n685), .ZN(G3) );
  NOR2_X1 U752 ( .A1(n704), .A2(n689), .ZN(n688) );
  XNOR2_X1 U753 ( .A(G104), .B(KEYINPUT113), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(G6) );
  NOR2_X1 U755 ( .A1(n706), .A2(n689), .ZN(n694) );
  XOR2_X1 U756 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n691) );
  XNOR2_X1 U757 ( .A(G107), .B(KEYINPUT114), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(KEYINPUT26), .B(n692), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n694), .B(n693), .ZN(G9) );
  XOR2_X1 U761 ( .A(n695), .B(G110), .Z(G12) );
  XOR2_X1 U762 ( .A(G128), .B(KEYINPUT29), .Z(n698) );
  NAND2_X1 U763 ( .A1(n701), .A2(n696), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(G30) );
  XNOR2_X1 U765 ( .A(G143), .B(n699), .ZN(G45) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(KEYINPUT116), .ZN(n703) );
  XNOR2_X1 U768 ( .A(G146), .B(n703), .ZN(G48) );
  NOR2_X1 U769 ( .A1(n707), .A2(n704), .ZN(n705) );
  XOR2_X1 U770 ( .A(G113), .B(n705), .Z(G15) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U772 ( .A(G116), .B(n708), .Z(G18) );
  XOR2_X1 U773 ( .A(G125), .B(KEYINPUT37), .Z(n709) );
  XNOR2_X1 U774 ( .A(n710), .B(n709), .ZN(G27) );
  XNOR2_X1 U775 ( .A(G134), .B(n711), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(KEYINPUT117), .ZN(G36) );
  INV_X1 U777 ( .A(n714), .ZN(n762) );
  NAND2_X1 U778 ( .A1(n762), .A2(n632), .ZN(n715) );
  XNOR2_X1 U779 ( .A(n715), .B(KEYINPUT88), .ZN(n718) );
  NAND2_X1 U780 ( .A1(n716), .A2(n632), .ZN(n717) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n719), .B(KEYINPUT85), .ZN(n722) );
  NAND2_X1 U783 ( .A1(n720), .A2(KEYINPUT2), .ZN(n721) );
  NAND2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n760) );
  NOR2_X1 U785 ( .A1(n723), .A2(n400), .ZN(n724) );
  XNOR2_X1 U786 ( .A(KEYINPUT50), .B(n724), .ZN(n732) );
  XOR2_X1 U787 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n728) );
  NAND2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U789 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U790 ( .A1(n729), .A2(n597), .ZN(n730) );
  XOR2_X1 U791 ( .A(KEYINPUT119), .B(n730), .Z(n731) );
  NOR2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U794 ( .A(KEYINPUT51), .B(n735), .ZN(n736) );
  NAND2_X1 U795 ( .A1(n736), .A2(n754), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U798 ( .A(n742), .B(KEYINPUT120), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U800 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U801 ( .A1(n755), .A2(n747), .ZN(n748) );
  NAND2_X1 U802 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U803 ( .A(KEYINPUT52), .B(n750), .Z(n751) );
  NOR2_X1 U804 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U805 ( .A(n753), .B(KEYINPUT121), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U808 ( .A1(G953), .A2(n758), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U810 ( .A(KEYINPUT53), .B(n761), .Z(G75) );
  NOR2_X1 U811 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U812 ( .A(n763), .B(KEYINPUT125), .ZN(n768) );
  NAND2_X1 U813 ( .A1(G224), .A2(G953), .ZN(n764) );
  XNOR2_X1 U814 ( .A(n764), .B(KEYINPUT124), .ZN(n765) );
  XNOR2_X1 U815 ( .A(KEYINPUT61), .B(n765), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n766), .A2(G898), .ZN(n767) );
  NAND2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n769), .B(KEYINPUT127), .ZN(n777) );
  XNOR2_X1 U819 ( .A(G101), .B(KEYINPUT126), .ZN(n771) );
  XNOR2_X1 U820 ( .A(n772), .B(n771), .ZN(n773) );
  XNOR2_X1 U821 ( .A(n770), .B(n773), .ZN(n775) );
  NOR2_X1 U822 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U823 ( .A(n777), .B(n776), .Z(G69) );
  XOR2_X1 U824 ( .A(n778), .B(G122), .Z(G24) );
  XNOR2_X1 U825 ( .A(G137), .B(n779), .ZN(G39) );
  XNOR2_X1 U826 ( .A(G131), .B(n780), .ZN(G33) );
endmodule

