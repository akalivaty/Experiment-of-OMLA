//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n224), .A2(new_n207), .A3(new_n225), .ZN(new_n226));
  NOR4_X1   g0026(.A1(new_n212), .A2(new_n222), .A3(new_n223), .A4(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n225), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n247), .A2(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G50), .A2(G58), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n207), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n246), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n246), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n206), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n256), .B(new_n260), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n270), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n279), .B2(G223), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n206), .A2(G274), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT68), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT68), .A2(G41), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(G226), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n267), .B(new_n269), .C1(new_n293), .C2(G200), .ZN(new_n294));
  OAI211_X1 g0094(.A(G190), .B(new_n292), .C1(new_n280), .C2(new_n282), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT72), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n294), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n289), .B1(G244), .B2(new_n291), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n203), .B2(new_n270), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n279), .B2(G238), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n306), .B2(new_n282), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n247), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(KEYINPUT70), .B2(new_n250), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(KEYINPUT70), .B2(new_n250), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(new_n248), .B1(new_n207), .B2(new_n273), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n246), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n261), .A2(G77), .A3(new_n263), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(G77), .C2(new_n257), .ZN(new_n318));
  OR3_X1    g0118(.A1(new_n308), .A2(new_n310), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n318), .B(new_n321), .C1(G179), .C2(new_n307), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n293), .A2(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n283), .A2(new_n325), .A3(new_n292), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n265), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n302), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT77), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n282), .A2(G232), .A3(new_n290), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT76), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n282), .A2(new_n290), .A3(new_n333), .A4(G232), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n289), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G33), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n337), .A2(new_n339), .A3(G226), .A4(G1698), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n337), .A2(new_n339), .A3(G223), .A4(new_n271), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n282), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n335), .A2(G179), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n320), .B1(new_n335), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n330), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n332), .A2(new_n334), .ZN(new_n349));
  INV_X1    g0149(.A(new_n289), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G169), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n335), .A2(G179), .A3(new_n345), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n270), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n337), .A2(new_n339), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n254), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n254), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G58), .A2(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(G20), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G159), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n251), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n357), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  INV_X1    g0170(.A(new_n246), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n359), .A2(new_n361), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(G68), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n357), .C1(new_n362), .C2(new_n368), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n311), .A2(new_n263), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n262), .A2(new_n378), .B1(new_n257), .B2(new_n311), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n355), .A2(new_n356), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n356), .B1(new_n355), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n351), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G190), .B2(new_n351), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n377), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n377), .A2(new_n387), .A3(KEYINPUT17), .A4(new_n380), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT78), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n270), .A2(G226), .A3(new_n271), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT73), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT73), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(G33), .A3(G97), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n344), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n289), .B1(G238), .B2(new_n291), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT74), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G169), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(G169), .A4(new_n411), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(G179), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n258), .A2(new_n254), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT12), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n254), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n273), .B2(new_n248), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT11), .A3(new_n246), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n261), .A2(G68), .A3(new_n263), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT11), .B1(new_n421), .B2(new_n246), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n309), .B1(new_n405), .B2(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n409), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n410), .A2(G200), .A3(new_n411), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n329), .A2(new_n394), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT5), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n285), .B2(new_n286), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n206), .A2(G45), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT5), .ZN(new_n441));
  AOI21_X1  g0241(.A(G41), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n436), .B(new_n438), .C1(new_n442), .C2(KEYINPUT84), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT84), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n444), .A2(new_n445), .A3(G41), .ZN(new_n446));
  OAI211_X1 g0246(.A(G270), .B(new_n282), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(KEYINPUT84), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n444), .B2(G41), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT68), .B(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n437), .B1(new_n450), .B2(new_n435), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n282), .A2(G274), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n449), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT88), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT88), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n447), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n270), .A2(G257), .A3(new_n271), .ZN(new_n458));
  INV_X1    g0258(.A(G303), .ZN(new_n459));
  INV_X1    g0259(.A(G264), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n458), .B1(new_n459), .B2(new_n270), .C1(new_n275), .C2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n455), .A2(new_n457), .B1(new_n344), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n257), .A2(new_n463), .A3(new_n225), .A4(new_n245), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n258), .A2(KEYINPUT89), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT89), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n257), .B2(G116), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n465), .A2(G116), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT91), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n471), .A2(KEYINPUT20), .B1(new_n207), .B2(G116), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n371), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT90), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n202), .A2(KEYINPUT80), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G97), .ZN(new_n477));
  AOI21_X1  g0277(.A(G33), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n207), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n480), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT80), .B(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(KEYINPUT90), .C1(new_n483), .C2(G33), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n473), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n470), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n481), .A2(new_n484), .ZN(new_n490));
  INV_X1    g0290(.A(new_n473), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n490), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT21), .B(G169), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT92), .B1(new_n462), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n461), .A2(new_n344), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n447), .A2(new_n456), .A3(new_n453), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n456), .B1(new_n447), .B2(new_n453), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n470), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n490), .A2(new_n491), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n487), .ZN(new_n501));
  INV_X1    g0301(.A(new_n492), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n320), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT92), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n498), .A2(new_n503), .A3(new_n504), .A4(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n503), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n489), .A2(new_n492), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n325), .B1(new_n461), .B2(new_n344), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n455), .A2(new_n457), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(G200), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n509), .C1(new_n309), .C2(new_n498), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n443), .A2(new_n446), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n337), .A2(new_n339), .A3(G244), .A4(new_n271), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n337), .A2(new_n339), .A3(G250), .A4(G1698), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n479), .A4(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n518), .A2(new_n452), .B1(new_n524), .B2(new_n344), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G257), .A3(new_n282), .ZN(new_n527));
  AOI21_X1  g0327(.A(G169), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n479), .B(new_n523), .C1(new_n519), .C2(new_n520), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n344), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n531), .A3(new_n325), .A4(new_n453), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n204), .A2(KEYINPUT81), .A3(new_n537), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n475), .A2(new_n477), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n543), .A2(new_n535), .A3(new_n203), .ZN(new_n544));
  OAI21_X1  g0344(.A(G20), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n251), .A2(new_n273), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(KEYINPUT82), .B1(G107), .B2(new_n372), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT82), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n371), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n258), .A2(new_n202), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n464), .B2(new_n202), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n534), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n535), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n538), .A2(new_n539), .A3(new_n536), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT81), .B1(new_n204), .B2(new_n537), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n543), .A2(new_n535), .A3(new_n203), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n207), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT82), .B1(new_n561), .B2(new_n546), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n372), .A2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n551), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n246), .ZN(new_n565));
  INV_X1    g0365(.A(new_n554), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n527), .A2(new_n453), .A3(new_n531), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n525), .A2(G190), .A3(new_n527), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n565), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n437), .A2(G250), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n344), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n337), .A2(new_n339), .A3(G244), .A4(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n270), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G116), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n574), .B1(new_n581), .B2(new_n344), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n320), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n325), .B(new_n574), .C1(new_n581), .C2(new_n344), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT86), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(G179), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n320), .C2(new_n582), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT19), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n207), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G87), .A2(G107), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n483), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n483), .B2(new_n248), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n270), .A2(new_n207), .A3(G68), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(KEYINPUT87), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n589), .A2(new_n207), .B1(new_n483), .B2(new_n591), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n601), .A3(new_n246), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n314), .A2(new_n258), .ZN(new_n603));
  INV_X1    g0403(.A(new_n314), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n465), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n585), .A2(new_n588), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n582), .A2(new_n309), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G200), .B2(new_n582), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n465), .A2(G87), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n603), .A4(new_n602), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n526), .A2(G264), .A3(new_n282), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n270), .A2(G250), .A3(new_n271), .ZN(new_n614));
  INV_X1    g0414(.A(G294), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n614), .C1(new_n336), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n344), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(new_n453), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(new_n617), .A3(G190), .A4(new_n453), .ZN(new_n620));
  OR3_X1    g0420(.A1(new_n257), .A2(KEYINPUT25), .A3(G107), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT25), .B1(new_n257), .B2(G107), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n203), .C2(new_n464), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT94), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n337), .A2(new_n339), .A3(new_n207), .A4(G87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT22), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT22), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n270), .A2(new_n628), .A3(new_n207), .A4(G87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT23), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n203), .A3(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT93), .ZN(new_n633));
  NAND2_X1  g0433(.A1(KEYINPUT23), .A2(G107), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n632), .A2(KEYINPUT93), .B1(new_n636), .B2(G20), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT24), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n630), .A2(new_n638), .A3(KEYINPUT24), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n246), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n619), .A2(new_n620), .A3(new_n625), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n625), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n612), .A2(new_n617), .A3(new_n325), .A4(new_n453), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n618), .A2(new_n320), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n607), .A2(new_n611), .A3(new_n644), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n571), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n434), .A2(new_n515), .A3(new_n517), .A4(new_n650), .ZN(G372));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(new_n606), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n583), .A2(new_n584), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n582), .A2(G200), .ZN(new_n655));
  AOI211_X1 g0455(.A(G190), .B(new_n574), .C1(new_n581), .C2(new_n344), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n602), .A2(new_n610), .A3(new_n603), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n653), .A2(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n652), .B1(new_n555), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT95), .B(new_n652), .C1(new_n555), .C2(new_n659), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n527), .A2(new_n453), .A3(new_n531), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n532), .B1(new_n664), .B2(G169), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n565), .B2(new_n566), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .A3(new_n611), .A4(new_n607), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n654), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n606), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n506), .A2(new_n514), .A3(new_n648), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n555), .A2(new_n570), .A3(new_n611), .A4(new_n644), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n434), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n390), .A2(new_n391), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT78), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n391), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n416), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n426), .B1(new_n683), .B2(new_n415), .ZN(new_n684));
  INV_X1    g0484(.A(new_n432), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n322), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n681), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n352), .A2(new_n353), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n381), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(new_n356), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n327), .B1(new_n691), .B2(new_n302), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n676), .A2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(G13), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n207), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n698), .A3(new_n207), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n492), .B2(new_n489), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n515), .A2(new_n517), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n515), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n648), .A2(new_n706), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n645), .A2(new_n706), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n644), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n648), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n648), .ZN(new_n717));
  NOR4_X1   g0517(.A1(new_n515), .A2(new_n717), .A3(new_n706), .A4(new_n714), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n712), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n210), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n450), .ZN(new_n722));
  INV_X1    g0522(.A(new_n224), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n592), .A2(G116), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G1), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n612), .A2(new_n617), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n664), .A2(new_n730), .A3(new_n510), .A4(new_n582), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n496), .A2(new_n497), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n582), .A2(G179), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(new_n618), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n498), .A3(new_n567), .ZN(new_n736));
  AND4_X1   g0536(.A1(new_n510), .A2(new_n582), .A3(new_n612), .A4(new_n617), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n513), .A2(new_n737), .A3(KEYINPUT30), .A4(new_n664), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n706), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n706), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n515), .A2(new_n650), .A3(new_n517), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(KEYINPUT31), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n733), .A2(new_n736), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n749), .A2(new_n738), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  AOI211_X1 g0554(.A(KEYINPUT29), .B(new_n706), .C1(new_n668), .C2(new_n674), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n672), .A2(new_n673), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n607), .A2(new_n611), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n652), .B1(new_n758), .B2(new_n555), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n666), .A2(KEYINPUT26), .A3(new_n611), .A4(new_n670), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n670), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n756), .B1(new_n762), .B2(new_n742), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT98), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n754), .A2(KEYINPUT98), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n728), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n694), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n206), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n722), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n711), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n709), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n210), .A2(new_n270), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n210), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n721), .A2(new_n270), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n288), .B2(new_n723), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n240), .A2(new_n288), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n225), .B1(G20), .B2(new_n320), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n774), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(new_n325), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G190), .A3(new_n385), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n207), .A2(G179), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n385), .A2(G190), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n793), .A2(new_n363), .B1(new_n796), .B2(new_n203), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n309), .A2(new_n385), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n797), .B1(G50), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT99), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G190), .A2(G200), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n792), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(new_n792), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n792), .A2(new_n795), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n801), .B1(new_n273), .B2(new_n806), .C1(new_n254), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n794), .A2(new_n803), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n367), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n798), .A2(new_n794), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n360), .B1(new_n817), .B2(G87), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n207), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n815), .B(new_n818), .C1(new_n202), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G326), .A2(new_n800), .B1(new_n817), .B2(G303), .ZN(new_n822));
  INV_X1    g0622(.A(new_n796), .ZN(new_n823));
  INV_X1    g0623(.A(new_n813), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n823), .A2(G283), .B1(new_n824), .B2(G329), .ZN(new_n825));
  INV_X1    g0625(.A(new_n793), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n270), .B1(new_n826), .B2(G322), .ZN(new_n827));
  INV_X1    g0627(.A(new_n820), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G294), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n822), .A2(new_n825), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(KEYINPUT33), .B(G317), .Z(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n811), .A2(new_n831), .B1(new_n832), .B2(new_n806), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n812), .A2(new_n821), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n788), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n791), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n787), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n709), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n776), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n323), .A2(new_n742), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n675), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n706), .B1(new_n668), .B2(new_n674), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n322), .A2(new_n706), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n318), .A2(new_n706), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n319), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n850), .B2(new_n322), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n846), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n754), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n774), .B1(new_n754), .B2(new_n852), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n851), .A2(new_n786), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n788), .A2(new_n785), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n774), .B1(G77), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n826), .A2(G143), .B1(new_n800), .B2(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n860), .B1(new_n367), .B2(new_n806), .C1(new_n811), .C2(new_n249), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT34), .Z(new_n862));
  AOI21_X1  g0662(.A(new_n360), .B1(new_n817), .B2(G50), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n828), .A2(G58), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n823), .A2(G68), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n824), .A2(G132), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n820), .A2(new_n202), .B1(new_n793), .B2(new_n615), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT102), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n800), .A2(G303), .B1(new_n824), .B2(G311), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n203), .B2(new_n816), .ZN(new_n871));
  INV_X1    g0671(.A(G87), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n796), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n871), .A2(new_n270), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G283), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n466), .B2(new_n806), .C1(new_n875), .C2(new_n811), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n862), .A2(new_n867), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n859), .B1(new_n877), .B2(new_n788), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n542), .A2(new_n544), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n225), .A2(new_n207), .A3(new_n466), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  OAI211_X1 g0687(.A(new_n723), .B(G77), .C1(new_n363), .C2(new_n254), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n259), .A2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n206), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n374), .A2(new_n369), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n892), .A2(new_n379), .ZN(new_n893));
  INV_X1    g0693(.A(new_n704), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n394), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n892), .A2(new_n379), .B1(new_n688), .B2(new_n894), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n388), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n704), .B(KEYINPUT105), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n381), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n388), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n355), .B2(new_n381), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n910), .B(new_n907), .C1(new_n394), .C2(new_n896), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n740), .A2(KEYINPUT107), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n739), .A2(new_n914), .A3(new_n706), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n745), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n739), .A2(new_n746), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n743), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n427), .A2(new_n706), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT103), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n433), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n428), .A2(new_n432), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(new_n851), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n912), .A2(new_n925), .A3(KEYINPUT40), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n428), .B2(new_n432), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n684), .A2(new_n685), .A3(new_n920), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n851), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n743), .A2(new_n917), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n916), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n377), .A2(new_n380), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n348), .A2(new_n354), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT18), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n355), .A2(new_n356), .A3(new_n381), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n679), .B2(new_n680), .ZN(new_n938));
  OAI211_X1 g0738(.A(KEYINPUT38), .B(new_n908), .C1(new_n938), .C2(new_n895), .ZN(new_n939));
  INV_X1    g0739(.A(new_n677), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n902), .B1(new_n690), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n689), .A2(new_n902), .A3(new_n388), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n903), .A2(new_n906), .B1(new_n942), .B2(new_n905), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n910), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n927), .B1(new_n932), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n926), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n434), .A2(new_n918), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(G330), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n844), .B1(new_n668), .B2(new_n674), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n924), .B1(new_n952), .B2(new_n848), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT104), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT104), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(new_n924), .C1(new_n952), .C2(new_n848), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n895), .B1(new_n681), .B2(new_n384), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n910), .B1(new_n957), .B2(new_n907), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n939), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n690), .A2(new_n901), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n945), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(KEYINPUT39), .A3(new_n939), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n428), .A2(new_n706), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n960), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n434), .B1(new_n755), .B2(new_n763), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n692), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n951), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n206), .B2(new_n771), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n951), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n891), .B1(new_n973), .B2(new_n974), .ZN(G367));
  NOR2_X1   g0775(.A1(new_n515), .A2(new_n706), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n715), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n706), .B1(new_n552), .B2(new_n554), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n555), .A2(new_n978), .A3(new_n570), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n666), .A2(new_n706), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT42), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n981), .B(KEYINPUT108), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n666), .B1(new_n985), .B2(new_n717), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n706), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n658), .A2(new_n706), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n670), .A2(new_n611), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n670), .B2(new_n988), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(KEYINPUT43), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT109), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT109), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n987), .A2(new_n995), .A3(new_n992), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n985), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n716), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT111), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n712), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n977), .A2(new_n1002), .A3(new_n981), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n719), .B2(new_n981), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT44), .B(new_n982), .C1(new_n718), .C2(new_n712), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1005), .A2(new_n1009), .A3(new_n716), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n716), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT110), .B1(new_n976), .B2(new_n715), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n711), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n710), .B(KEYINPUT110), .C1(new_n715), .C2(new_n976), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n718), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n718), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1013), .A2(new_n1019), .B1(new_n767), .B2(new_n768), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n722), .B(KEYINPUT41), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n1001), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n772), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1020), .A2(new_n1001), .A3(new_n1021), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1000), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n781), .A2(new_n235), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n789), .B1(new_n210), .B2(new_n314), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n774), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n816), .A2(new_n1029), .A3(new_n466), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n360), .B1(new_n813), .B2(new_n1031), .C1(new_n483), .C2(new_n796), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G107), .C2(new_n828), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n826), .A2(G303), .B1(new_n800), .B2(G311), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(KEYINPUT112), .B2(new_n1034), .C1(new_n615), .C2(new_n811), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n816), .B2(new_n466), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1034), .A2(KEYINPUT112), .B1(KEYINPUT113), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(KEYINPUT113), .B2(new_n1036), .C1(new_n875), .C2(new_n806), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n793), .A2(new_n249), .B1(new_n816), .B2(new_n363), .ZN(new_n1039));
  INV_X1    g0839(.A(G143), .ZN(new_n1040));
  INV_X1    g0840(.A(G137), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n799), .A2(new_n1040), .B1(new_n813), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n820), .A2(new_n254), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n270), .B1(new_n796), .B2(new_n273), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n259), .B2(new_n806), .C1(new_n367), .C2(new_n811), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1035), .A2(new_n1038), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT47), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1028), .B1(new_n1049), .B2(new_n788), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n840), .B2(new_n990), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1025), .A2(new_n1051), .ZN(G387));
  XNOR2_X1  g0852(.A(new_n725), .B(KEYINPUT115), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n288), .B1(new_n254), .B2(new_n273), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n247), .A2(G50), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1053), .B(new_n1057), .C1(new_n1056), .C2(new_n1055), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n780), .C1(new_n288), .C2(new_n231), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(G107), .B2(new_n210), .C1(new_n725), .C2(new_n777), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n722), .B(new_n773), .C1(new_n1060), .C2(new_n789), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n811), .A2(new_n247), .B1(new_n254), .B2(new_n806), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n793), .A2(new_n259), .B1(new_n813), .B2(new_n249), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n799), .A2(new_n367), .B1(new_n796), .B2(new_n202), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n270), .B1(new_n816), .B2(new_n273), .C1(new_n820), .C2(new_n314), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n826), .A2(G317), .B1(new_n800), .B2(G322), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n459), .B2(new_n806), .C1(new_n811), .C2(new_n832), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n828), .A2(G283), .B1(new_n817), .B2(G294), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT49), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g0875(.A(G326), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n360), .B1(new_n813), .B2(new_n1076), .C1(new_n466), .C2(new_n796), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1074), .B2(KEYINPUT116), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1066), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1061), .B1(new_n715), .B2(new_n840), .C1(new_n1079), .C2(new_n837), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1019), .A2(new_n769), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n722), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1019), .A2(new_n769), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1080), .B1(new_n772), .B2(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n722), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1081), .B1(new_n767), .B2(new_n768), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n1013), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1082), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n780), .A2(new_n243), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n790), .B1(new_n721), .B2(new_n543), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n722), .B(new_n773), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n793), .A2(new_n832), .B1(new_n799), .B2(new_n1031), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT52), .Z(new_n1096));
  OAI22_X1  g0896(.A1(new_n811), .A2(new_n459), .B1(new_n615), .B2(new_n806), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G283), .A2(new_n817), .B1(new_n824), .B2(G322), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(new_n360), .C1(new_n203), .C2(new_n796), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n820), .A2(new_n466), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n806), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n311), .B1(G77), .B2(new_n828), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n259), .B2(new_n811), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT117), .Z(new_n1105));
  OAI22_X1  g0905(.A1(new_n793), .A2(new_n367), .B1(new_n799), .B2(new_n249), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI22_X1  g0907(.A1(new_n816), .A2(new_n254), .B1(new_n813), .B2(new_n1040), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1107), .A2(new_n360), .A3(new_n873), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1101), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1094), .B1(new_n837), .B2(new_n1110), .C1(new_n985), .C2(new_n840), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1013), .B2(new_n773), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1090), .A2(new_n1091), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1091), .B1(new_n1090), .B2(new_n1113), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G390));
  INV_X1    g0917(.A(new_n966), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n964), .A2(new_n965), .B1(new_n953), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT119), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n966), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n945), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n928), .A2(new_n929), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n850), .A2(new_n322), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n762), .A2(new_n742), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n848), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT120), .B1(new_n1119), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n706), .B1(new_n674), .B2(new_n761), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n848), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n945), .B(new_n1123), .C1(new_n1134), .C2(new_n1125), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT39), .B1(new_n939), .B2(new_n944), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n912), .B2(KEYINPUT39), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n846), .A2(new_n1128), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n966), .B1(new_n1138), .B2(new_n924), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1132), .B(new_n1135), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n918), .A2(new_n924), .A3(G330), .A4(new_n851), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1131), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT121), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n753), .A2(G330), .A3(new_n851), .A4(new_n924), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n1135), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1131), .A2(new_n1140), .A3(KEYINPUT121), .A4(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n434), .A2(G330), .A3(new_n918), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n969), .A2(new_n1150), .A3(new_n692), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT122), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n969), .A2(new_n1150), .A3(KEYINPUT122), .A4(new_n692), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(G330), .B(new_n851), .C1(new_n744), .C2(new_n752), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1125), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1141), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n918), .A2(G330), .A3(new_n851), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1125), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1159), .A2(new_n1138), .B1(new_n1146), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1156), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1149), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1155), .A2(new_n1163), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n722), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1137), .A2(new_n786), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1102), .A2(new_n1172), .B1(G159), .B2(new_n828), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1041), .B2(new_n811), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT123), .Z(new_n1175));
  AOI22_X1  g0975(.A1(new_n826), .A2(G132), .B1(new_n824), .B2(G125), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n799), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n249), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT53), .B1(new_n816), .B2(new_n249), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n270), .C1(new_n259), .C2(new_n796), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1175), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n360), .B1(new_n816), .B2(new_n872), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n793), .A2(new_n466), .B1(new_n799), .B2(new_n875), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G77), .C2(new_n828), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n203), .B2(new_n811), .C1(new_n483), .C2(new_n806), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n865), .B1(new_n615), .B2(new_n813), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT124), .Z(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n788), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n774), .C1(new_n311), .C2(new_n858), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1170), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n773), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1169), .A2(new_n1194), .ZN(G378));
  AOI22_X1  g0995(.A1(G125), .A2(new_n800), .B1(new_n817), .B2(new_n1172), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1177), .B2(new_n793), .ZN(new_n1197));
  INV_X1    g0997(.A(G132), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n811), .A2(new_n1198), .B1(new_n1041), .B2(new_n806), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(G150), .C2(new_n828), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n824), .A2(G124), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n823), .C2(G159), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n811), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1207), .A2(G97), .B1(new_n604), .B2(new_n1102), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n796), .A2(new_n363), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n793), .A2(new_n203), .B1(new_n813), .B2(new_n875), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G116), .C2(new_n800), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n360), .B(new_n287), .C1(new_n816), .C2(new_n273), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(new_n1043), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n259), .B1(G33), .B2(G41), .C1(new_n270), .C2(new_n450), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1218));
  AND4_X1   g1018(.A1(new_n1206), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n774), .B1(G50), .B2(new_n858), .C1(new_n1219), .C2(new_n837), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n302), .A2(new_n328), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n894), .A2(new_n265), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT55), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1221), .B(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(KEYINPUT125), .B(KEYINPUT56), .Z(new_n1225));
  XNOR2_X1  g1025(.A(new_n1224), .B(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1226), .B2(new_n785), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT126), .Z(new_n1228));
  OAI21_X1  g1028(.A(G330), .B1(new_n926), .B2(new_n946), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n961), .B1(new_n1137), .B2(new_n966), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n960), .ZN(new_n1231));
  INV_X1    g1031(.A(G330), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n945), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT40), .B1(new_n1233), .B2(new_n925), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n932), .A2(new_n927), .A3(new_n959), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n968), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1226), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1231), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1231), .B2(new_n1237), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1228), .B1(new_n1241), .B2(new_n773), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1168), .A2(new_n1156), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1239), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n722), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1243), .B2(new_n1241), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1242), .B1(new_n1247), .B2(new_n1248), .ZN(G375));
  INV_X1    g1049(.A(new_n1021), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1155), .A2(new_n1163), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1165), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n774), .B1(G68), .B2(new_n858), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n793), .A2(new_n875), .B1(new_n813), .B2(new_n459), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n811), .A2(new_n466), .B1(new_n203), .B2(new_n806), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n799), .A2(new_n615), .B1(new_n816), .B2(new_n202), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n360), .B1(new_n796), .B2(new_n273), .C1(new_n820), .C2(new_n314), .ZN(new_n1257));
  OR4_X1    g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1207), .A2(new_n1172), .B1(G150), .B2(new_n1102), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n826), .A2(G137), .B1(new_n824), .B2(G128), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G132), .A2(new_n800), .B1(new_n817), .B2(G159), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n360), .B(new_n1209), .C1(G50), .C2(new_n828), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1253), .B1(new_n1267), .B2(new_n788), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n924), .B2(new_n786), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1163), .B2(new_n772), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1252), .A2(new_n1271), .ZN(G381));
  NOR4_X1   g1072(.A1(G393), .A2(G396), .A3(G381), .A4(G384), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1116), .A2(new_n1273), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G387), .A2(new_n1274), .A3(G378), .A4(G375), .ZN(G407));
  OAI22_X1  g1075(.A1(new_n1149), .A2(new_n772), .B1(new_n1170), .B2(new_n1191), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1086), .B1(new_n1149), .B2(new_n1165), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1168), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n705), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(G387), .A2(new_n1116), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(G393), .B(new_n842), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1025), .B(new_n1051), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1242), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1243), .A2(new_n1250), .A3(new_n1241), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1227), .B1(new_n1241), .B2(new_n773), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1278), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1279), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1280), .A2(G2897), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1155), .A2(new_n1163), .A3(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n722), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1251), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n879), .B1(new_n1301), .B2(new_n1270), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1301), .A2(new_n879), .A3(new_n1270), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1297), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1302), .A3(new_n1296), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1295), .B2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1280), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1288), .A2(new_n1310), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1315), .A2(new_n1318), .A3(new_n1312), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1315), .B2(new_n1308), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1315), .B2(new_n1312), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1323), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1278), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1313), .A3(new_n1289), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1313), .B1(new_n1325), .B2(new_n1289), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1288), .ZN(G402));
endmodule


