//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(new_n457), .B1(G567), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(new_n457), .B2(new_n456), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT65), .Z(G319));
  AND2_X1   g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G125), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n466), .B(G2105), .C1(new_n472), .C2(new_n461), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(G160));
  NAND2_X1  g054(.A1(new_n476), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND2_X1  g061(.A1(new_n481), .A2(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n464), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n471), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n464), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n476), .A2(new_n496), .A3(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT69), .B(new_n499), .C1(new_n500), .C2(KEYINPUT68), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n500), .B2(KEYINPUT69), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n509), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT7), .Z(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n506), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n510), .A2(new_n511), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n499), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT69), .B1(new_n500), .B2(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n527), .B2(new_n501), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n512), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g107(.A(KEYINPUT70), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(G52), .A2(new_n534), .B1(new_n528), .B2(G90), .ZN(new_n538));
  AND2_X1   g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n506), .B2(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n540), .B2(new_n508), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n527), .B2(new_n501), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n542), .B(G651), .C1(new_n544), .C2(new_n539), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n534), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n528), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n506), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n508), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT72), .B1(new_n528), .B2(G91), .ZN(new_n562));
  AND4_X1   g137(.A1(KEYINPUT72), .A2(new_n506), .A3(G91), .A4(new_n515), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n506), .B2(G65), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n508), .B1(new_n568), .B2(KEYINPUT73), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n527), .B2(new_n501), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n572), .B2(new_n567), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(KEYINPUT74), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT74), .B1(new_n569), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n538), .A2(new_n541), .A3(new_n579), .A4(new_n545), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n528), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n513), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n528), .A2(G86), .B1(G48), .B2(new_n513), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n508), .B2(new_n589), .ZN(G305));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT70), .B1(new_n515), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n533), .ZN(new_n593));
  OAI21_X1  g168(.A(G47), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n506), .A2(G85), .A3(new_n515), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n506), .A2(G60), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n508), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n527), .B2(new_n501), .ZN(new_n602));
  INV_X1    g177(.A(new_n598), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n604), .A2(KEYINPUT76), .A3(new_n594), .A4(new_n595), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(new_n534), .A2(G54), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT77), .B(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n527), .B2(new_n501), .ZN(new_n609));
  AND2_X1   g184(.A1(G79), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(KEYINPUT10), .B1(new_n528), .B2(G92), .ZN(new_n612));
  AND4_X1   g187(.A1(KEYINPUT10), .A2(new_n506), .A3(G92), .A4(new_n515), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n607), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n581), .B2(G868), .ZN(G284));
  XOR2_X1   g191(.A(G284), .B(KEYINPUT78), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n568), .A2(KEYINPUT73), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n620), .A2(new_n573), .A3(G651), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n564), .B1(new_n623), .B2(new_n574), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(G868), .B2(new_n624), .ZN(G297));
  OAI21_X1  g200(.A(new_n619), .B1(G868), .B2(new_n624), .ZN(G280));
  INV_X1    g201(.A(new_n614), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g208(.A1(new_n469), .A2(G2105), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n462), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(new_n640));
  INV_X1    g215(.A(new_n637), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n481), .A2(G123), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT81), .Z(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(G111), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G2105), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(G135), .B2(new_n476), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n641), .A2(G2100), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n640), .B(new_n650), .C1(new_n642), .C2(new_n649), .ZN(G156));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n638), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n642), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(new_n696), .B(new_n695), .S(new_n688), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1981), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n685), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n704), .A3(new_n685), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n683), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(new_n683), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n709), .A2(new_n710), .A3(new_n705), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  XOR2_X1   g288(.A(KEYINPUT85), .B(G16), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT88), .Z(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(G6), .A2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(G305), .B2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n723), .A2(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n719), .A2(new_n726), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT90), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n715), .A2(G24), .ZN(new_n737));
  XNOR2_X1  g312(.A(G290), .B(KEYINPUT86), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n715), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1986), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n733), .A2(new_n734), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G25), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n476), .A2(G131), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G119), .ZN(new_n745));
  OR2_X1    g320(.A1(G95), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n742), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  XOR2_X1   g326(.A(new_n750), .B(new_n751), .Z(new_n752));
  OR4_X1    g327(.A1(new_n736), .A2(new_n740), .A3(new_n741), .A4(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n462), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n464), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n476), .A2(G139), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n742), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n742), .B2(G33), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G35), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G162), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT29), .B(G2090), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT30), .B(G28), .ZN(new_n772));
  OR2_X1    g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n772), .A2(new_n742), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n649), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n742), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n769), .B2(new_n770), .ZN(new_n778));
  NOR2_X1   g353(.A1(G164), .A2(new_n742), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G27), .B2(new_n742), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n771), .B(new_n784), .C1(new_n767), .C2(new_n766), .ZN(new_n785));
  NAND2_X1  g360(.A1(G168), .A2(G16), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(KEYINPUT95), .C1(G16), .C2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT95), .B2(new_n786), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G1966), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n742), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n476), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n481), .A2(G128), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G29), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(KEYINPUT92), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n728), .A2(G5), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G171), .B2(new_n728), .ZN(new_n804));
  INV_X1    g379(.A(G1961), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n785), .A2(new_n789), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n788), .A2(G1966), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT96), .ZN(new_n809));
  OR2_X1    g384(.A1(KEYINPUT24), .A2(G34), .ZN(new_n810));
  NAND2_X1  g385(.A1(KEYINPUT24), .A2(G34), .ZN(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G160), .B2(G29), .ZN(new_n813));
  INV_X1    g388(.A(G2084), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G4), .A2(G16), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n627), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1348), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n715), .A2(G19), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n554), .B2(new_n715), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1341), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n742), .A2(G32), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n634), .A2(new_n824), .A3(G105), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT93), .ZN(new_n827));
  AOI22_X1  g402(.A1(G141), .A2(new_n476), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n481), .A2(G129), .ZN(new_n829));
  NAND3_X1  g404(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT26), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT26), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n828), .A2(KEYINPUT94), .A3(new_n829), .A4(new_n833), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n823), .B1(new_n838), .B2(new_n742), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT27), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1996), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n809), .A2(new_n815), .A3(new_n822), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n714), .A2(G20), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G299), .B2(G16), .ZN(new_n846));
  INV_X1    g421(.A(G1956), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n807), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n755), .A2(new_n756), .A3(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  AND2_X1   g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n506), .B2(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n854), .B2(new_n508), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n527), .B2(new_n501), .ZN(new_n857));
  OAI211_X1 g432(.A(KEYINPUT98), .B(G651), .C1(new_n857), .C2(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(G55), .A2(new_n534), .B1(new_n528), .B2(G93), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n627), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n550), .A2(KEYINPUT99), .A3(new_n553), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  AOI22_X1  g442(.A1(G43), .A2(new_n534), .B1(new_n528), .B2(G81), .ZN(new_n868));
  INV_X1    g443(.A(G56), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n527), .B2(new_n501), .ZN(new_n870));
  INV_X1    g445(.A(new_n552), .ZN(new_n871));
  OAI21_X1  g446(.A(G651), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n867), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n861), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT99), .B1(new_n550), .B2(new_n553), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n867), .A3(new_n872), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n875), .A2(new_n859), .A3(new_n860), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n865), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n882));
  INV_X1    g457(.A(G860), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n863), .B1(new_n881), .B2(new_n884), .ZN(G145));
  AND2_X1   g460(.A1(G160), .A2(G162), .ZN(new_n886));
  NOR2_X1   g461(.A1(G160), .A2(G162), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(new_n649), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n886), .A2(new_n887), .A3(new_n776), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n476), .A2(G142), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n481), .A2(G130), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n464), .A2(G118), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n636), .B(new_n896), .ZN(new_n897));
  MUX2_X1   g472(.A(KEYINPUT102), .B(KEYINPUT101), .S(new_n764), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n497), .A2(new_n495), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n488), .A2(new_n489), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n481), .B2(G126), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n898), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n838), .B(new_n796), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(new_n748), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n898), .A2(new_n902), .ZN(new_n909));
  INV_X1    g484(.A(new_n897), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n748), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n906), .A2(new_n908), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n911), .A2(new_n906), .B1(new_n908), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n891), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n906), .A2(new_n911), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n913), .C1(new_n890), .C2(new_n889), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n924));
  NAND2_X1  g499(.A1(G166), .A2(G305), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n589), .A2(new_n508), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(new_n588), .C1(new_n509), .C2(new_n518), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n600), .A2(new_n605), .A3(new_n722), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n722), .B1(new_n600), .B2(new_n605), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n924), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n928), .B1(new_n933), .B2(KEYINPUT103), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n878), .B(new_n630), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n623), .A2(new_n574), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n627), .B1(new_n940), .B2(new_n565), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n564), .B(new_n614), .C1(new_n623), .C2(new_n574), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(G299), .A2(new_n614), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n624), .A2(new_n627), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n944), .B1(new_n939), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n938), .B1(new_n951), .B2(KEYINPUT104), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(KEYINPUT104), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n952), .B(new_n953), .ZN(new_n954));
  MUX2_X1   g529(.A(new_n861), .B(new_n954), .S(G868), .Z(G295));
  MUX2_X1   g530(.A(new_n861), .B(new_n954), .S(G868), .Z(G331));
  NAND2_X1  g531(.A1(new_n581), .A2(G168), .ZN(new_n957));
  NAND2_X1  g532(.A1(G286), .A2(new_n546), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n878), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G286), .B1(new_n578), .B2(new_n580), .ZN(new_n960));
  AND2_X1   g535(.A1(G286), .A2(new_n546), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n877), .B(new_n874), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n943), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n959), .A2(new_n962), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n936), .B(new_n963), .C1(new_n964), .C2(new_n950), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n921), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n964), .B2(new_n950), .ZN(new_n968));
  INV_X1    g543(.A(new_n936), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n968), .A2(KEYINPUT105), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT105), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n966), .B(new_n967), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(KEYINPUT105), .A3(new_n969), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n967), .A4(new_n966), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n967), .B1(new_n966), .B2(new_n974), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n973), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n984));
  INV_X1    g559(.A(new_n966), .ZN(new_n985));
  INV_X1    g560(.A(new_n974), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n967), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  MUX2_X1   g563(.A(new_n983), .B(new_n988), .S(KEYINPUT44), .Z(G397));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n476), .A2(G137), .ZN(new_n991));
  INV_X1    g566(.A(new_n475), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(G40), .A3(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n990), .B(new_n993), .C1(new_n465), .C2(new_n473), .ZN(new_n994));
  INV_X1    g569(.A(new_n993), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT107), .B1(new_n474), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(G164), .B2(G1384), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT124), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1000), .B(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g581(.A(new_n838), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n796), .B(new_n801), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1005), .B(new_n1010), .C1(new_n1003), .C2(new_n1002), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(new_n838), .B2(new_n1001), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n748), .B(new_n751), .Z(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1006), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1000), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1012), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n749), .A2(new_n751), .ZN(new_n1024));
  OAI22_X1  g599(.A1(new_n1015), .A2(new_n1024), .B1(G2067), .B2(new_n796), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1006), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n999), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n997), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n474), .A2(new_n995), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n990), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n474), .A2(KEYINPUT107), .A3(new_n995), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n902), .A2(new_n1040), .A3(new_n1032), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n902), .A2(new_n1032), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1039), .A2(new_n814), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1035), .A2(new_n1044), .A3(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1030), .B1(new_n1049), .B2(G168), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(G8), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G286), .A2(G8), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1027), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1028), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT120), .B1(new_n1057), .B2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT62), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1052), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1057), .A2(KEYINPUT120), .A3(new_n1054), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1048), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT119), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1067));
  OAI21_X1  g642(.A(G168), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1029), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1061), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT55), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n902), .B2(new_n1032), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n998), .B(G1384), .C1(new_n899), .C2(new_n901), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1971), .B1(new_n1039), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1043), .B(new_n1079), .C1(new_n994), .C2(new_n996), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1041), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2090), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1074), .B1(new_n1085), .B2(new_n1028), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1042), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n994), .B2(new_n996), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT110), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1092), .B1(G1976), .B2(new_n722), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n926), .A2(new_n701), .A3(new_n588), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n589), .A2(new_n508), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n513), .A2(G48), .ZN(new_n1103));
  INV_X1    g678(.A(G86), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n516), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n701), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1100), .A2(new_n1101), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1107), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT49), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1111), .B2(new_n1099), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1093), .A2(new_n1095), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1074), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1043), .B(new_n1041), .C1(new_n994), .C2(new_n996), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1078), .A2(KEYINPUT109), .B1(G2090), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1078), .A2(KEYINPUT109), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1116), .B(G8), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1092), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1091), .B1(new_n1088), .B2(G8), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1121), .A2(new_n1122), .B1(new_n1094), .B2(G288), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT52), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1086), .A2(new_n1115), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1039), .A2(new_n1077), .A3(new_n781), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1117), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1039), .A2(KEYINPUT115), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n805), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1062), .A2(new_n1072), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G288), .A2(G1976), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1096), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1114), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1124), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1120), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1140), .B(KEYINPUT112), .C1(new_n1120), .C2(new_n1143), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1057), .A2(G168), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1125), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1149), .B(new_n1150), .C1(new_n1152), .C2(new_n1074), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n1120), .A3(new_n1124), .A4(new_n1115), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1135), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n847), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT56), .B(G2072), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1039), .A2(new_n1077), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n624), .A2(KEYINPUT114), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n624), .B2(KEYINPUT114), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1158), .A2(new_n1160), .A3(new_n1164), .A4(new_n1163), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1157), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  INV_X1    g744(.A(G1348), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1129), .A2(new_n1130), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1039), .A2(new_n801), .A3(new_n1087), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n627), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n614), .A3(new_n1172), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1169), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n997), .A2(new_n1034), .A3(G1996), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT58), .B(G1341), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1039), .B2(new_n1087), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n554), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n554), .B(new_n1181), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n627), .A2(new_n1169), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1183), .B(new_n1184), .C1(new_n1173), .C2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1168), .A2(new_n1176), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1161), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1158), .A2(KEYINPUT116), .A3(new_n1160), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1165), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(KEYINPUT61), .A3(new_n1167), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1174), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1187), .A2(new_n1192), .B1(new_n1193), .B2(new_n1167), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1070), .A2(new_n1125), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT54), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT53), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT53), .B(new_n781), .C1(new_n463), .C2(new_n464), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n993), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1126), .A2(new_n1197), .B1(new_n1077), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1131), .A2(new_n1200), .A3(G301), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1196), .B1(new_n1132), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(KEYINPUT121), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1204), .B(new_n1196), .C1(new_n1132), .C2(new_n1201), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1127), .A2(G301), .A3(new_n1131), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1131), .A2(new_n1200), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(G171), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1207), .A2(new_n1209), .A3(KEYINPUT54), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(KEYINPUT122), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1207), .A2(new_n1209), .A3(new_n1212), .A4(KEYINPUT54), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1195), .A2(new_n1206), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT123), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1194), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1195), .A2(new_n1206), .A3(KEYINPUT123), .A4(new_n1214), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1156), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(G290), .B(new_n703), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1017), .B1(new_n1018), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1026), .B1(new_n1219), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g797(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1224));
  XNOR2_X1  g798(.A(new_n1224), .B(KEYINPUT126), .ZN(new_n1225));
  NAND3_X1  g799(.A1(new_n712), .A2(new_n1225), .A3(new_n922), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n981), .B1(new_n972), .B2(KEYINPUT106), .ZN(new_n1227));
  AOI211_X1 g801(.A(KEYINPUT127), .B(new_n1226), .C1(new_n1227), .C2(new_n980), .ZN(new_n1228));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1229));
  INV_X1    g803(.A(new_n1226), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1229), .B1(new_n983), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g805(.A1(new_n1228), .A2(new_n1231), .ZN(G308));
  NAND2_X1  g806(.A1(new_n983), .A2(new_n1230), .ZN(G225));
endmodule


