

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799;

  XNOR2_X1 U368 ( .A(n571), .B(KEYINPUT108), .ZN(n759) );
  NAND2_X1 U369 ( .A1(n620), .A2(n610), .ZN(n744) );
  XNOR2_X1 U370 ( .A(G131), .B(G140), .ZN(n543) );
  XNOR2_X1 U371 ( .A(G113), .B(G122), .ZN(n545) );
  INV_X2 U372 ( .A(KEYINPUT64), .ZN(n659) );
  AND2_X2 U373 ( .A1(n600), .A2(n425), .ZN(n424) );
  NAND2_X2 U374 ( .A1(n397), .A2(n418), .ZN(n444) );
  XNOR2_X2 U375 ( .A(n346), .B(n591), .ZN(n436) );
  NAND2_X2 U376 ( .A1(n366), .A2(n365), .ZN(n346) );
  XNOR2_X1 U377 ( .A(G134), .B(G107), .ZN(n523) );
  NAND2_X1 U378 ( .A1(G234), .A2(G237), .ZN(n480) );
  INV_X1 U379 ( .A(G237), .ZN(n501) );
  INV_X1 U380 ( .A(G902), .ZN(n457) );
  INV_X2 U381 ( .A(G140), .ZN(n676) );
  XNOR2_X2 U382 ( .A(n615), .B(n614), .ZN(n644) );
  NAND2_X2 U383 ( .A1(n563), .A2(n763), .ZN(n405) );
  XNOR2_X2 U384 ( .A(n504), .B(KEYINPUT77), .ZN(n563) );
  NOR2_X2 U385 ( .A1(n589), .A2(n744), .ZN(n437) );
  AND2_X2 U386 ( .A1(n435), .A2(n432), .ZN(n431) );
  XOR2_X1 U387 ( .A(KEYINPUT123), .B(n703), .Z(n704) );
  NAND2_X2 U388 ( .A1(n670), .A2(n668), .ZN(n571) );
  NOR2_X2 U389 ( .A1(G953), .A2(G237), .ZN(n490) );
  NAND2_X1 U390 ( .A1(n439), .A2(n652), .ZN(n438) );
  OR2_X1 U391 ( .A1(n599), .A2(n422), .ZN(n636) );
  XNOR2_X1 U392 ( .A(n606), .B(KEYINPUT0), .ZN(n613) );
  AND2_X1 U393 ( .A1(n570), .A2(n564), .ZN(n609) );
  XNOR2_X1 U394 ( .A(n522), .B(n521), .ZN(n594) );
  XNOR2_X1 U395 ( .A(n688), .B(G116), .ZN(n524) );
  XNOR2_X1 U396 ( .A(G119), .B(G110), .ZN(n466) );
  NAND2_X1 U397 ( .A1(n408), .A2(n410), .ZN(n417) );
  NAND2_X1 U398 ( .A1(n347), .A2(n656), .ZN(n741) );
  NAND2_X1 U399 ( .A1(n430), .A2(n434), .ZN(n429) );
  AND2_X1 U400 ( .A1(n355), .A2(n367), .ZN(n365) );
  NAND2_X1 U401 ( .A1(n419), .A2(n352), .ZN(n418) );
  AND2_X1 U402 ( .A1(n398), .A2(n441), .ZN(n397) );
  XNOR2_X1 U403 ( .A(n561), .B(n389), .ZN(n402) );
  XNOR2_X1 U404 ( .A(n390), .B(KEYINPUT113), .ZN(n368) );
  OR2_X1 U405 ( .A1(n636), .A2(n428), .ZN(n357) );
  NAND2_X1 U406 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U407 ( .A(n679), .B(n680), .ZN(n681) );
  BUF_X1 U408 ( .A(n594), .Z(n404) );
  NAND2_X1 U409 ( .A1(n594), .A2(n762), .ZN(n568) );
  XNOR2_X1 U410 ( .A(n660), .B(KEYINPUT59), .ZN(n661) );
  XNOR2_X1 U411 ( .A(n713), .B(n714), .ZN(n715) );
  XOR2_X1 U412 ( .A(KEYINPUT122), .B(n707), .Z(n708) );
  XNOR2_X1 U413 ( .A(n370), .B(n720), .ZN(n721) );
  XNOR2_X1 U414 ( .A(n510), .B(KEYINPUT10), .ZN(n787) );
  XOR2_X2 U415 ( .A(KEYINPUT107), .B(KEYINPUT9), .Z(n526) );
  XNOR2_X1 U416 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n461) );
  INV_X2 U417 ( .A(G122), .ZN(n688) );
  XNOR2_X2 U418 ( .A(G110), .B(G107), .ZN(n450) );
  XNOR2_X2 U419 ( .A(KEYINPUT15), .B(G902), .ZN(n517) );
  XNOR2_X1 U420 ( .A(KEYINPUT89), .B(KEYINPUT46), .ZN(n562) );
  XNOR2_X2 U421 ( .A(G119), .B(G101), .ZN(n494) );
  XNOR2_X1 U422 ( .A(KEYINPUT7), .B(KEYINPUT106), .ZN(n525) );
  INV_X1 U423 ( .A(KEYINPUT8), .ZN(n459) );
  XNOR2_X1 U424 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n462) );
  INV_X4 U425 ( .A(G953), .ZN(n792) );
  BUF_X2 U426 ( .A(n719), .Z(n711) );
  INV_X1 U427 ( .A(n409), .ZN(n347) );
  AND2_X2 U428 ( .A1(n790), .A2(n348), .ZN(n409) );
  XNOR2_X2 U429 ( .A(n438), .B(n653), .ZN(n348) );
  XNOR2_X1 U430 ( .A(n438), .B(n653), .ZN(n693) );
  BUF_X1 U431 ( .A(n555), .Z(n349) );
  OR2_X2 U432 ( .A1(n396), .A2(n426), .ZN(n423) );
  XNOR2_X2 U433 ( .A(n403), .B(n659), .ZN(n719) );
  OR2_X2 U434 ( .A1(n679), .A2(G902), .ZN(n361) );
  NAND2_X1 U435 ( .A1(n414), .A2(n412), .ZN(n411) );
  NAND2_X1 U436 ( .A1(n517), .A2(n415), .ZN(n414) );
  NAND2_X1 U437 ( .A1(n654), .A2(n413), .ZN(n412) );
  NAND2_X1 U438 ( .A1(KEYINPUT2), .A2(n415), .ZN(n413) );
  NAND2_X1 U439 ( .A1(n402), .A2(n387), .ZN(n399) );
  OR2_X1 U440 ( .A1(n402), .A2(n387), .ZN(n401) );
  XNOR2_X1 U441 ( .A(G113), .B(KEYINPUT70), .ZN(n495) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n509) );
  OR2_X2 U443 ( .A1(n370), .A2(n654), .ZN(n522) );
  BUF_X1 U444 ( .A(n619), .Z(n751) );
  XNOR2_X1 U445 ( .A(n393), .B(n359), .ZN(n392) );
  INV_X1 U446 ( .A(KEYINPUT65), .ZN(n415) );
  XNOR2_X1 U447 ( .A(n400), .B(n580), .ZN(n367) );
  NAND2_X1 U448 ( .A1(n354), .A2(n579), .ZN(n400) );
  XOR2_X1 U449 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n473) );
  AND2_X1 U450 ( .A1(n656), .A2(KEYINPUT65), .ZN(n416) );
  INV_X1 U451 ( .A(KEYINPUT87), .ZN(n434) );
  AND2_X1 U452 ( .A1(n433), .A2(n675), .ZN(n432) );
  NAND2_X1 U453 ( .A1(n677), .A2(n434), .ZN(n433) );
  NAND2_X1 U454 ( .A1(n422), .A2(KEYINPUT110), .ZN(n421) );
  XNOR2_X1 U455 ( .A(G137), .B(KEYINPUT5), .ZN(n488) );
  XOR2_X1 U456 ( .A(G116), .B(KEYINPUT102), .Z(n489) );
  XNOR2_X1 U457 ( .A(G101), .B(KEYINPUT78), .ZN(n452) );
  XNOR2_X1 U458 ( .A(G134), .B(G131), .ZN(n448) );
  INV_X1 U459 ( .A(KEYINPUT30), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n619), .B(KEYINPUT6), .ZN(n645) );
  XNOR2_X1 U461 ( .A(n516), .B(n690), .ZN(n370) );
  NOR2_X1 U462 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U463 ( .A(n608), .ZN(n442) );
  AND2_X1 U464 ( .A1(n613), .A2(KEYINPUT34), .ZN(n443) );
  INV_X1 U465 ( .A(n748), .ZN(n394) );
  INV_X1 U466 ( .A(KEYINPUT42), .ZN(n389) );
  INV_X1 U467 ( .A(n621), .ZN(n395) );
  AND2_X1 U468 ( .A1(n640), .A2(n428), .ZN(n641) );
  XNOR2_X1 U469 ( .A(n402), .B(n388), .ZN(G39) );
  INV_X1 U470 ( .A(G137), .ZN(n388) );
  INV_X1 U471 ( .A(n445), .ZN(n422) );
  XOR2_X1 U472 ( .A(n500), .B(G472), .Z(n350) );
  XOR2_X1 U473 ( .A(n475), .B(n474), .Z(n351) );
  AND2_X1 U474 ( .A1(n371), .A2(n607), .ZN(n352) );
  XOR2_X1 U475 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n353) );
  AND2_X1 U476 ( .A1(n577), .A2(n667), .ZN(n354) );
  AND2_X1 U477 ( .A1(n399), .A2(n739), .ZN(n355) );
  AND2_X1 U478 ( .A1(n445), .A2(n426), .ZN(n356) );
  AND2_X1 U479 ( .A1(n597), .A2(KEYINPUT87), .ZN(n358) );
  XOR2_X1 U480 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n359) );
  INV_X1 U481 ( .A(n562), .ZN(n387) );
  AND2_X1 U482 ( .A1(n654), .A2(n415), .ZN(n360) );
  INV_X1 U483 ( .A(n645), .ZN(n600) );
  XNOR2_X2 U484 ( .A(n361), .B(n350), .ZN(n619) );
  NAND2_X1 U485 ( .A1(n363), .A2(n362), .ZN(n366) );
  NAND2_X1 U486 ( .A1(n686), .A2(n401), .ZN(n362) );
  NAND2_X1 U487 ( .A1(n385), .A2(n562), .ZN(n363) );
  AND2_X2 U488 ( .A1(n368), .A2(n369), .ZN(n671) );
  NAND2_X1 U489 ( .A1(n756), .A2(n368), .ZN(n561) );
  NAND2_X1 U490 ( .A1(n369), .A2(n605), .ZN(n606) );
  XNOR2_X2 U491 ( .A(n568), .B(KEYINPUT19), .ZN(n369) );
  INV_X1 U492 ( .A(n613), .ZN(n371) );
  XNOR2_X2 U493 ( .A(n403), .B(n659), .ZN(n372) );
  BUF_X1 U494 ( .A(n515), .Z(n373) );
  INV_X1 U495 ( .A(n599), .ZN(n374) );
  BUF_X1 U496 ( .A(n759), .Z(n375) );
  INV_X1 U497 ( .A(n396), .ZN(n599) );
  AND2_X2 U498 ( .A1(n423), .A2(n421), .ZN(n420) );
  XNOR2_X1 U499 ( .A(n589), .B(n353), .ZN(n396) );
  INV_X1 U500 ( .A(n600), .ZN(n376) );
  BUF_X1 U501 ( .A(n589), .Z(n377) );
  NOR2_X1 U502 ( .A1(n655), .A2(n656), .ZN(n657) );
  NAND2_X1 U503 ( .A1(n409), .A2(n360), .ZN(n408) );
  NAND2_X1 U504 ( .A1(n790), .A2(n381), .ZN(n378) );
  NAND2_X1 U505 ( .A1(n378), .A2(n379), .ZN(n410) );
  OR2_X1 U506 ( .A1(n380), .A2(n416), .ZN(n379) );
  INV_X1 U507 ( .A(n411), .ZN(n380) );
  AND2_X1 U508 ( .A1(n693), .A2(n411), .ZN(n381) );
  XNOR2_X1 U509 ( .A(n784), .B(G146), .ZN(n382) );
  XNOR2_X1 U510 ( .A(n784), .B(G146), .ZN(n499) );
  XNOR2_X1 U511 ( .A(n407), .B(n406), .ZN(n502) );
  XNOR2_X2 U512 ( .A(G146), .B(G125), .ZN(n510) );
  XNOR2_X2 U513 ( .A(n383), .B(n384), .ZN(n589) );
  NOR2_X1 U514 ( .A1(n712), .A2(G902), .ZN(n383) );
  XOR2_X1 U515 ( .A(n458), .B(KEYINPUT68), .Z(n384) );
  XNOR2_X2 U516 ( .A(n658), .B(KEYINPUT76), .ZN(n742) );
  NAND2_X2 U517 ( .A1(n417), .A2(n742), .ZN(n403) );
  INV_X1 U518 ( .A(n686), .ZN(n385) );
  XNOR2_X2 U519 ( .A(n386), .B(KEYINPUT40), .ZN(n686) );
  NAND2_X2 U520 ( .A1(n555), .A2(n554), .ZN(n386) );
  INV_X1 U521 ( .A(n377), .ZN(n391) );
  NAND2_X1 U522 ( .A1(n427), .A2(n619), .ZN(n393) );
  NAND2_X1 U523 ( .A1(n356), .A2(n396), .ZN(n425) );
  NAND2_X1 U524 ( .A1(n599), .A2(n394), .ZN(n646) );
  NAND2_X1 U525 ( .A1(n395), .A2(n599), .ZN(n622) );
  NAND2_X1 U526 ( .A1(n590), .A2(n374), .ZN(n739) );
  NAND2_X1 U527 ( .A1(n758), .A2(KEYINPUT34), .ZN(n398) );
  XNOR2_X2 U528 ( .A(n602), .B(n601), .ZN(n758) );
  INV_X1 U529 ( .A(n581), .ZN(n427) );
  NAND2_X2 U530 ( .A1(n431), .A2(n429), .ZN(n655) );
  XNOR2_X1 U531 ( .A(n437), .B(KEYINPUT101), .ZN(n639) );
  XNOR2_X2 U532 ( .A(n405), .B(KEYINPUT39), .ZN(n555) );
  NAND2_X1 U533 ( .A1(n619), .A2(n762), .ZN(n407) );
  INV_X1 U534 ( .A(n620), .ZN(n748) );
  XNOR2_X2 U535 ( .A(n476), .B(n351), .ZN(n620) );
  INV_X1 U536 ( .A(n758), .ZN(n419) );
  NAND2_X2 U537 ( .A1(n424), .A2(n420), .ZN(n602) );
  INV_X1 U538 ( .A(KEYINPUT110), .ZN(n426) );
  INV_X1 U539 ( .A(n751), .ZN(n428) );
  NAND2_X1 U540 ( .A1(n436), .A2(n358), .ZN(n435) );
  INV_X1 U541 ( .A(n436), .ZN(n430) );
  INV_X1 U542 ( .A(n349), .ZN(n598) );
  XNOR2_X1 U543 ( .A(n440), .B(n651), .ZN(n439) );
  NAND2_X1 U544 ( .A1(n650), .A2(n649), .ZN(n440) );
  XNOR2_X2 U545 ( .A(n444), .B(KEYINPUT35), .ZN(n689) );
  INV_X1 U546 ( .A(n744), .ZN(n445) );
  BUF_X1 U547 ( .A(n758), .Z(n779) );
  NOR2_X1 U548 ( .A1(n617), .A2(n616), .ZN(n446) );
  AND2_X1 U549 ( .A1(n685), .A2(n678), .ZN(n624) );
  INV_X1 U550 ( .A(KEYINPUT48), .ZN(n591) );
  INV_X1 U551 ( .A(KEYINPUT71), .ZN(n626) );
  XNOR2_X1 U552 ( .A(n627), .B(n626), .ZN(n629) );
  XNOR2_X1 U553 ( .A(n382), .B(n498), .ZN(n679) );
  INV_X1 U554 ( .A(KEYINPUT60), .ZN(n665) );
  XNOR2_X2 U555 ( .A(G128), .B(KEYINPUT80), .ZN(n447) );
  XNOR2_X2 U556 ( .A(n447), .B(G143), .ZN(n532) );
  XNOR2_X2 U557 ( .A(n532), .B(KEYINPUT4), .ZN(n515) );
  XNOR2_X1 U558 ( .A(n448), .B(KEYINPUT67), .ZN(n449) );
  XNOR2_X2 U559 ( .A(n515), .B(n449), .ZN(n784) );
  XNOR2_X1 U560 ( .A(n450), .B(G104), .ZN(n505) );
  NAND2_X1 U561 ( .A1(n792), .A2(G227), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U563 ( .A(n505), .B(n453), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n676), .B(G137), .ZN(n467) );
  INV_X1 U565 ( .A(n467), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n454), .B(KEYINPUT95), .ZN(n786) );
  XOR2_X1 U567 ( .A(n455), .B(n786), .Z(n456) );
  XNOR2_X1 U568 ( .A(n499), .B(n456), .ZN(n712) );
  XNOR2_X1 U569 ( .A(KEYINPUT69), .B(G469), .ZN(n458) );
  NAND2_X1 U570 ( .A1(n792), .A2(G234), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n460), .B(n459), .ZN(n529) );
  NAND2_X1 U572 ( .A1(n529), .A2(G221), .ZN(n464) );
  XNOR2_X1 U573 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U574 ( .A(n464), .B(n463), .ZN(n471) );
  XNOR2_X2 U575 ( .A(G128), .B(KEYINPUT23), .ZN(n465) );
  XNOR2_X1 U576 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U578 ( .A(n469), .B(n787), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n470), .B(n471), .ZN(n703) );
  OR2_X2 U580 ( .A1(n703), .A2(G902), .ZN(n476) );
  NAND2_X1 U581 ( .A1(G234), .A2(n517), .ZN(n472) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n477) );
  NAND2_X1 U583 ( .A1(n477), .A2(G217), .ZN(n475) );
  XNOR2_X1 U584 ( .A(KEYINPUT100), .B(KEYINPUT25), .ZN(n474) );
  NAND2_X1 U585 ( .A1(n477), .A2(G221), .ZN(n479) );
  INV_X1 U586 ( .A(KEYINPUT21), .ZN(n478) );
  XNOR2_X1 U587 ( .A(n479), .B(n478), .ZN(n610) );
  XNOR2_X1 U588 ( .A(n480), .B(KEYINPUT14), .ZN(n772) );
  INV_X1 U589 ( .A(G952), .ZN(n663) );
  NAND2_X1 U590 ( .A1(n792), .A2(n663), .ZN(n482) );
  OR2_X1 U591 ( .A1(n792), .A2(G902), .ZN(n481) );
  AND2_X1 U592 ( .A1(n482), .A2(n481), .ZN(n483) );
  AND2_X1 U593 ( .A1(n772), .A2(n483), .ZN(n604) );
  NAND2_X1 U594 ( .A1(G953), .A2(G900), .ZN(n484) );
  NAND2_X1 U595 ( .A1(n604), .A2(n484), .ZN(n486) );
  INV_X1 U596 ( .A(KEYINPUT82), .ZN(n485) );
  XNOR2_X1 U597 ( .A(n486), .B(n485), .ZN(n556) );
  INV_X1 U598 ( .A(n556), .ZN(n487) );
  NOR2_X1 U599 ( .A1(n639), .A2(n487), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n489), .B(n488), .ZN(n493) );
  INV_X1 U601 ( .A(n490), .ZN(n491) );
  XNOR2_X1 U602 ( .A(KEYINPUT75), .B(n491), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n538), .A2(G210), .ZN(n492) );
  XNOR2_X1 U604 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n494), .B(KEYINPUT3), .ZN(n496) );
  XNOR2_X1 U606 ( .A(n496), .B(n495), .ZN(n507) );
  XNOR2_X1 U607 ( .A(n497), .B(n507), .ZN(n498) );
  INV_X1 U608 ( .A(KEYINPUT72), .ZN(n500) );
  NAND2_X1 U609 ( .A1(n501), .A2(n457), .ZN(n518) );
  NAND2_X1 U610 ( .A1(n518), .A2(G214), .ZN(n762) );
  NAND2_X1 U611 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n524), .B(KEYINPUT16), .ZN(n506) );
  XNOR2_X1 U613 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U614 ( .A(n508), .B(n507), .ZN(n690) );
  XNOR2_X1 U615 ( .A(n510), .B(n509), .ZN(n513) );
  NAND2_X1 U616 ( .A1(n792), .A2(G224), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n511), .B(KEYINPUT93), .ZN(n512) );
  XNOR2_X1 U618 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U619 ( .A(n373), .B(n514), .ZN(n516) );
  INV_X1 U620 ( .A(n517), .ZN(n654) );
  NAND2_X1 U621 ( .A1(n518), .A2(G210), .ZN(n520) );
  XNOR2_X1 U622 ( .A(KEYINPUT81), .B(KEYINPUT94), .ZN(n519) );
  XNOR2_X1 U623 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U624 ( .A(n404), .B(KEYINPUT38), .ZN(n760) );
  INV_X1 U625 ( .A(n760), .ZN(n763) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n528) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U628 ( .A(n528), .B(n527), .Z(n531) );
  NAND2_X1 U629 ( .A1(G217), .A2(n529), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n531), .B(n530), .ZN(n535) );
  BUF_X1 U631 ( .A(n532), .Z(n533) );
  INV_X1 U632 ( .A(n533), .ZN(n534) );
  XNOR2_X1 U633 ( .A(n535), .B(n534), .ZN(n707) );
  NAND2_X1 U634 ( .A1(n707), .A2(n457), .ZN(n537) );
  INV_X1 U635 ( .A(G478), .ZN(n536) );
  XNOR2_X1 U636 ( .A(n537), .B(n536), .ZN(n570) );
  INV_X1 U637 ( .A(n570), .ZN(n565) );
  NAND2_X1 U638 ( .A1(n538), .A2(G214), .ZN(n540) );
  XNOR2_X1 U639 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U641 ( .A(n787), .B(n541), .ZN(n549) );
  INV_X1 U642 ( .A(G143), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n542), .B(G104), .ZN(n544) );
  XNOR2_X1 U644 ( .A(n544), .B(n543), .ZN(n547) );
  XNOR2_X1 U645 ( .A(n545), .B(KEYINPUT104), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U647 ( .A(n549), .B(n548), .ZN(n660) );
  OR2_X1 U648 ( .A1(n660), .A2(G902), .ZN(n553) );
  XNOR2_X1 U649 ( .A(G475), .B(KEYINPUT13), .ZN(n551) );
  INV_X1 U650 ( .A(KEYINPUT105), .ZN(n550) );
  XNOR2_X1 U651 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U652 ( .A(n553), .B(n552), .ZN(n564) );
  OR2_X1 U653 ( .A1(n565), .A2(n564), .ZN(n668) );
  INV_X1 U654 ( .A(n668), .ZN(n554) );
  AND2_X1 U655 ( .A1(n556), .A2(n610), .ZN(n557) );
  NAND2_X1 U656 ( .A1(n748), .A2(n557), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n609), .A2(n762), .ZN(n558) );
  OR2_X1 U658 ( .A1(n760), .A2(n558), .ZN(n560) );
  XNOR2_X1 U659 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n559) );
  XNOR2_X1 U660 ( .A(n560), .B(n559), .ZN(n756) );
  BUF_X1 U661 ( .A(n563), .Z(n567) );
  INV_X1 U662 ( .A(n564), .ZN(n569) );
  AND2_X1 U663 ( .A1(n565), .A2(n569), .ZN(n608) );
  AND2_X1 U664 ( .A1(n404), .A2(n608), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n667) );
  OR2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n670) );
  INV_X1 U667 ( .A(KEYINPUT84), .ZN(n572) );
  NOR2_X1 U668 ( .A1(n572), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U669 ( .A1(n759), .A2(n573), .ZN(n575) );
  OR2_X1 U670 ( .A1(n759), .A2(KEYINPUT84), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n671), .A2(n576), .ZN(n577) );
  NAND2_X1 U673 ( .A1(n671), .A2(n375), .ZN(n578) );
  NAND2_X1 U674 ( .A1(n578), .A2(KEYINPUT47), .ZN(n579) );
  INV_X1 U675 ( .A(KEYINPUT74), .ZN(n580) );
  OR2_X1 U676 ( .A1(n645), .A2(n581), .ZN(n582) );
  XNOR2_X1 U677 ( .A(n582), .B(KEYINPUT111), .ZN(n585) );
  INV_X1 U678 ( .A(n762), .ZN(n583) );
  NOR2_X1 U679 ( .A1(n668), .A2(n583), .ZN(n584) );
  AND2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n592) );
  NAND2_X1 U681 ( .A1(n592), .A2(n404), .ZN(n588) );
  XNOR2_X1 U682 ( .A(KEYINPUT36), .B(KEYINPUT92), .ZN(n586) );
  XNOR2_X1 U683 ( .A(n586), .B(KEYINPUT115), .ZN(n587) );
  XNOR2_X1 U684 ( .A(n588), .B(n587), .ZN(n590) );
  NAND2_X1 U685 ( .A1(n592), .A2(n599), .ZN(n593) );
  XNOR2_X1 U686 ( .A(n593), .B(KEYINPUT43), .ZN(n596) );
  INV_X1 U687 ( .A(n404), .ZN(n595) );
  AND2_X1 U688 ( .A1(n596), .A2(n595), .ZN(n677) );
  INV_X1 U689 ( .A(n677), .ZN(n597) );
  OR2_X1 U690 ( .A1(n598), .A2(n670), .ZN(n675) );
  XNOR2_X2 U691 ( .A(n655), .B(KEYINPUT85), .ZN(n790) );
  INV_X1 U692 ( .A(KEYINPUT33), .ZN(n601) );
  NAND2_X1 U693 ( .A1(G953), .A2(G898), .ZN(n603) );
  AND2_X1 U694 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U695 ( .A(KEYINPUT34), .ZN(n607) );
  INV_X1 U696 ( .A(n689), .ZN(n625) );
  INV_X1 U697 ( .A(n609), .ZN(n764) );
  INV_X1 U698 ( .A(n610), .ZN(n747) );
  NOR2_X1 U699 ( .A1(n764), .A2(n747), .ZN(n611) );
  XNOR2_X1 U700 ( .A(n611), .B(KEYINPUT109), .ZN(n612) );
  OR2_X2 U701 ( .A1(n613), .A2(n612), .ZN(n615) );
  XNOR2_X1 U702 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n614) );
  XNOR2_X1 U703 ( .A(n376), .B(KEYINPUT79), .ZN(n617) );
  OR2_X1 U704 ( .A1(n599), .A2(n620), .ZN(n616) );
  NAND2_X1 U705 ( .A1(n644), .A2(n446), .ZN(n618) );
  XNOR2_X2 U706 ( .A(n618), .B(KEYINPUT32), .ZN(n685) );
  INV_X1 U707 ( .A(n644), .ZN(n623) );
  OR2_X1 U708 ( .A1(n751), .A2(n620), .ZN(n621) );
  OR2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n678) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n627) );
  INV_X1 U711 ( .A(KEYINPUT44), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n633) );
  AND2_X1 U713 ( .A1(n626), .A2(KEYINPUT44), .ZN(n630) );
  AND2_X1 U714 ( .A1(n678), .A2(n630), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n685), .A2(n631), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n652) );
  NAND2_X1 U717 ( .A1(n689), .A2(KEYINPUT44), .ZN(n635) );
  INV_X1 U718 ( .A(KEYINPUT91), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n635), .B(n634), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n357), .A2(n613), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n637) );
  XNOR2_X1 U722 ( .A(n638), .B(n637), .ZN(n735) );
  INV_X1 U723 ( .A(n639), .ZN(n640) );
  AND2_X1 U724 ( .A1(n641), .A2(n371), .ZN(n728) );
  OR2_X1 U725 ( .A1(n735), .A2(n728), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n375), .B(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n646), .A2(n600), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n644), .A2(n647), .ZN(n674) );
  AND2_X1 U730 ( .A1(n648), .A2(n674), .ZN(n649) );
  INV_X1 U731 ( .A(KEYINPUT90), .ZN(n651) );
  XNOR2_X1 U732 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n653) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n348), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n372), .A2(G475), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n663), .A2(G953), .ZN(n723) );
  NAND2_X1 U738 ( .A1(n664), .A2(n723), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(G60) );
  XNOR2_X1 U740 ( .A(n667), .B(G143), .ZN(G45) );
  NAND2_X1 U741 ( .A1(n671), .A2(n554), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(G146), .ZN(G48) );
  INV_X1 U743 ( .A(n670), .ZN(n734) );
  NAND2_X1 U744 ( .A1(n671), .A2(n734), .ZN(n673) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G30) );
  XNOR2_X1 U747 ( .A(n674), .B(G101), .ZN(G3) );
  XNOR2_X1 U748 ( .A(n675), .B(G134), .ZN(G36) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(G42) );
  XNOR2_X1 U750 ( .A(n678), .B(G110), .ZN(G12) );
  NAND2_X1 U751 ( .A1(n719), .A2(G472), .ZN(n682) );
  XOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT62), .Z(n680) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n683), .A2(n723), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n684), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U756 ( .A(n685), .B(G119), .ZN(G21) );
  BUF_X1 U757 ( .A(n686), .Z(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(G131), .ZN(G33) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(G24) );
  INV_X1 U760 ( .A(n690), .ZN(n692) );
  NOR2_X1 U761 ( .A1(G898), .A2(n792), .ZN(n691) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n702) );
  INV_X1 U763 ( .A(n348), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n694), .A2(G953), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G224), .A2(G953), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n695), .B(KEYINPUT61), .ZN(n696) );
  XNOR2_X1 U767 ( .A(KEYINPUT124), .B(n696), .ZN(n697) );
  NAND2_X1 U768 ( .A1(n697), .A2(G898), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT125), .ZN(n699) );
  NOR2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U771 ( .A(n702), .B(n701), .Z(G69) );
  NAND2_X1 U772 ( .A1(n711), .A2(G217), .ZN(n705) );
  XNOR2_X1 U773 ( .A(n705), .B(n704), .ZN(n706) );
  INV_X1 U774 ( .A(n723), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n706), .A2(n717), .ZN(G66) );
  NAND2_X1 U776 ( .A1(n711), .A2(G478), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U778 ( .A1(n710), .A2(n717), .ZN(G63) );
  NAND2_X1 U779 ( .A1(n711), .A2(G469), .ZN(n716) );
  BUF_X1 U780 ( .A(n712), .Z(n713) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n714) );
  XNOR2_X1 U782 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n372), .A2(G210), .ZN(n722) );
  XNOR2_X1 U785 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n720) );
  XNOR2_X1 U786 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n726) );
  XOR2_X1 U788 ( .A(KEYINPUT88), .B(KEYINPUT56), .Z(n725) );
  XNOR2_X1 U789 ( .A(n726), .B(n725), .ZN(G51) );
  NAND2_X1 U790 ( .A1(n728), .A2(n554), .ZN(n727) );
  XNOR2_X1 U791 ( .A(n727), .B(G104), .ZN(G6) );
  XOR2_X1 U792 ( .A(KEYINPUT26), .B(KEYINPUT117), .Z(n730) );
  NAND2_X1 U793 ( .A1(n728), .A2(n734), .ZN(n729) );
  XNOR2_X1 U794 ( .A(n730), .B(n729), .ZN(n732) );
  XOR2_X1 U795 ( .A(G107), .B(KEYINPUT27), .Z(n731) );
  XNOR2_X1 U796 ( .A(n732), .B(n731), .ZN(G9) );
  NAND2_X1 U797 ( .A1(n735), .A2(n554), .ZN(n733) );
  XNOR2_X1 U798 ( .A(n733), .B(G113), .ZN(G15) );
  NAND2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U800 ( .A(n736), .B(KEYINPUT118), .ZN(n737) );
  XNOR2_X1 U801 ( .A(G116), .B(n737), .ZN(G18) );
  XNOR2_X1 U802 ( .A(KEYINPUT37), .B(KEYINPUT119), .ZN(n738) );
  XNOR2_X1 U803 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U804 ( .A(G125), .B(n740), .ZN(G27) );
  XOR2_X1 U805 ( .A(KEYINPUT83), .B(n741), .Z(n743) );
  NAND2_X1 U806 ( .A1(n743), .A2(n742), .ZN(n777) );
  XOR2_X1 U807 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n746) );
  NAND2_X1 U808 ( .A1(n599), .A2(n744), .ZN(n745) );
  XOR2_X1 U809 ( .A(n746), .B(n745), .Z(n753) );
  NAND2_X1 U810 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U811 ( .A(n749), .B(KEYINPUT49), .ZN(n750) );
  NOR2_X1 U812 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U813 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U814 ( .A1(n754), .A2(n357), .ZN(n755) );
  XNOR2_X1 U815 ( .A(KEYINPUT51), .B(n755), .ZN(n757) );
  INV_X1 U816 ( .A(n756), .ZN(n778) );
  NOR2_X1 U817 ( .A1(n757), .A2(n778), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n375), .A2(n762), .ZN(n761) );
  NOR2_X1 U819 ( .A1(n761), .A2(n760), .ZN(n767) );
  NOR2_X1 U820 ( .A1(n763), .A2(n762), .ZN(n765) );
  NOR2_X1 U821 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U822 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U823 ( .A1(n779), .A2(n768), .ZN(n769) );
  NOR2_X1 U824 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U825 ( .A(KEYINPUT52), .B(n771), .ZN(n774) );
  NAND2_X1 U826 ( .A1(G952), .A2(n772), .ZN(n773) );
  NOR2_X1 U827 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U828 ( .A1(G953), .A2(n775), .ZN(n776) );
  NAND2_X1 U829 ( .A1(n777), .A2(n776), .ZN(n782) );
  NOR2_X1 U830 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U831 ( .A(KEYINPUT121), .B(n780), .Z(n781) );
  NOR2_X1 U832 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U833 ( .A(KEYINPUT53), .B(n783), .ZN(G75) );
  BUF_X1 U834 ( .A(n784), .Z(n785) );
  XOR2_X1 U835 ( .A(KEYINPUT126), .B(n786), .Z(n788) );
  XNOR2_X1 U836 ( .A(n788), .B(n787), .ZN(n789) );
  XNOR2_X1 U837 ( .A(n785), .B(n789), .ZN(n794) );
  BUF_X1 U838 ( .A(n790), .Z(n791) );
  XOR2_X1 U839 ( .A(n794), .B(n791), .Z(n793) );
  NAND2_X1 U840 ( .A1(n793), .A2(n792), .ZN(n799) );
  XNOR2_X1 U841 ( .A(G227), .B(n794), .ZN(n795) );
  NAND2_X1 U842 ( .A1(n795), .A2(G900), .ZN(n796) );
  XOR2_X1 U843 ( .A(KEYINPUT127), .B(n796), .Z(n797) );
  NAND2_X1 U844 ( .A1(G953), .A2(n797), .ZN(n798) );
  NAND2_X1 U845 ( .A1(n799), .A2(n798), .ZN(G72) );
endmodule

