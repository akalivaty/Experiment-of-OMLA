//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n208), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  AND4_X1   g017(.A1(new_n210), .A2(new_n211), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n216), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT95), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(KEYINPUT95), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT96), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n209), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n225), .B2(new_n209), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n220), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n209), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT96), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n219), .B1(new_n233), .B2(new_n227), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT103), .ZN(new_n238));
  AND2_X1   g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(KEYINPUT103), .C1(KEYINPUT102), .C2(KEYINPUT7), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  INV_X1    g047(.A(G92gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(KEYINPUT8), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT102), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n241), .A2(new_n253), .A3(new_n243), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G99gat), .B(G106gat), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n246), .A2(new_n258), .A3(new_n250), .A4(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n237), .A2(new_n260), .B1(KEYINPUT41), .B2(new_n202), .ZN(new_n261));
  XNOR2_X1  g060(.A(G134gat), .B(G162gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n230), .A2(new_n259), .A3(new_n257), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n261), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n206), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n205), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G71gat), .A2(G78gat), .ZN(new_n273));
  OR2_X1    g072(.A1(G71gat), .A2(G78gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT9), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G57gat), .B(G64gat), .Z(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT101), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT101), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(KEYINPUT9), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n274), .A2(new_n273), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT100), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n274), .B(new_n273), .C1(new_n285), .C2(new_n275), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT100), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n280), .B(new_n281), .C1(new_n284), .C2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT21), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(KEYINPUT21), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT16), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(G1gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G1gat), .B2(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(G8gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n294), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n295), .B1(new_n294), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G231gat), .A3(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n302), .B2(new_n303), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n305), .B2(new_n307), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n293), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n314), .ZN(new_n316));
  INV_X1    g115(.A(new_n293), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n272), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT104), .ZN(new_n321));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G204gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n241), .A2(new_n253), .A3(new_n243), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n253), .B1(new_n241), .B2(new_n243), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n258), .B1(new_n330), .B2(new_n250), .ZN(new_n331));
  INV_X1    g130(.A(new_n259), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n289), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n286), .B(new_n287), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n280), .A2(new_n281), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n257), .A2(new_n334), .A3(new_n335), .A4(new_n259), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(KEYINPUT105), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT105), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n290), .A2(new_n338), .A3(new_n259), .A4(new_n257), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT106), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT106), .ZN(new_n346));
  AOI211_X1 g145(.A(new_n346), .B(KEYINPUT10), .C1(new_n337), .C2(new_n339), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n336), .A2(new_n344), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT107), .ZN(new_n350));
  INV_X1    g149(.A(new_n341), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n340), .A2(new_n344), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(new_n348), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT106), .A3(new_n344), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT107), .B1(new_n357), .B2(new_n341), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n327), .B(new_n343), .C1(new_n352), .C2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n326), .B(KEYINPUT108), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n349), .A2(new_n351), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n342), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT109), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(KEYINPUT109), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n321), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(G169gat), .B2(G176gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT24), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT64), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(G183gat), .B2(G190gat), .ZN(new_n376));
  INV_X1    g175(.A(G190gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n295), .A2(new_n377), .A3(KEYINPUT64), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  INV_X1    g179(.A(G169gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n323), .A3(KEYINPUT23), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT65), .ZN(new_n383));
  AND4_X1   g182(.A1(new_n372), .A2(new_n379), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n380), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT66), .ZN(new_n386));
  OR2_X1    g185(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n374), .B1(new_n389), .B2(G190gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n371), .A3(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n371), .A2(new_n384), .B1(new_n391), .B2(KEYINPUT25), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT28), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(KEYINPUT27), .A3(new_n388), .ZN(new_n395));
  OR2_X1    g194(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n397), .B2(new_n377), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT68), .B(G190gat), .C1(new_n395), .C2(new_n396), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT27), .B(G183gat), .Z(new_n401));
  OAI21_X1  g200(.A(KEYINPUT28), .B1(new_n401), .B2(G190gat), .ZN(new_n402));
  OR3_X1    g201(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n380), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n400), .A2(new_n373), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT69), .Z(new_n409));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(KEYINPUT70), .Z(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n411), .B2(KEYINPUT1), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT71), .B(G120gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G113gat), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n414), .A2(KEYINPUT72), .ZN(new_n415));
  INV_X1    g214(.A(G113gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G120gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n415), .A2(new_n418), .A3(new_n419), .A4(new_n408), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT73), .B1(new_n407), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n421), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n412), .A2(new_n420), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n392), .A2(new_n424), .A3(new_n425), .A4(new_n406), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n427), .B2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n434), .A2(new_n435), .B1(KEYINPUT32), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT75), .B(G71gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n441), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT33), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT32), .B(new_n446), .C1(new_n434), .C2(new_n435), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n432), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n432), .A3(new_n447), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT36), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g255(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n457));
  INV_X1    g256(.A(G218gat), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n456), .B(new_n457), .C1(new_n309), .C2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G197gat), .B(G204gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G211gat), .B(G218gat), .Z(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n461), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT79), .ZN(new_n466));
  XOR2_X1   g265(.A(G141gat), .B(G148gat), .Z(new_n467));
  INV_X1    g266(.A(G155gat), .ZN(new_n468));
  INV_X1    g267(.A(G162gat), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT2), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G155gat), .B(G162gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n465), .B2(KEYINPUT29), .ZN(new_n480));
  INV_X1    g279(.A(new_n473), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n478), .B(KEYINPUT85), .ZN(new_n487));
  INV_X1    g286(.A(new_n462), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n476), .B1(new_n461), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n462), .B1(new_n459), .B2(new_n460), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n474), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G22gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n486), .A2(G22gat), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G50gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n496), .B(new_n497), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n421), .A2(new_n481), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n421), .A2(new_n481), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n424), .A2(new_n473), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n510), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT84), .A3(new_n509), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(KEYINPUT5), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n481), .A2(KEYINPUT3), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n421), .A3(new_n475), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n521), .A2(new_n508), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT5), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT0), .B(G57gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G85gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G1gat), .B(G29gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT89), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n526), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n537), .A2(new_n509), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n509), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(KEYINPUT40), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(KEYINPUT40), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  NAND2_X1  g345(.A1(G226gat), .A2(G233gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT80), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n407), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n407), .B2(new_n476), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n466), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n466), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT29), .B1(new_n392), .B2(new_n406), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n549), .B(new_n553), .C1(new_n548), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(KEYINPUT81), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n551), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n553), .A4(new_n549), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G8gat), .B(G36gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G64gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n249), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT30), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT82), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n556), .A2(new_n559), .A3(new_n563), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n560), .A2(KEYINPUT82), .A3(KEYINPUT30), .A4(new_n564), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n567), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n536), .B(new_n546), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n578));
  INV_X1    g377(.A(new_n533), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n528), .B1(new_n519), .B2(new_n525), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n536), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT6), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT6), .A4(new_n579), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n564), .B1(new_n560), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n556), .A2(KEYINPUT37), .A3(new_n559), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n586), .B1(new_n587), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n552), .A2(new_n555), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT37), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n598), .A3(new_n589), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n596), .A2(KEYINPUT94), .B1(KEYINPUT92), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n594), .A2(new_n600), .A3(new_n568), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n507), .B1(new_n577), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT83), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n604), .A2(new_n605), .B1(new_n569), .B2(new_n568), .ZN(new_n606));
  INV_X1    g405(.A(new_n580), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT6), .B1(new_n607), .B2(new_n533), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n533), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n582), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n606), .B(new_n610), .C1(new_n605), .C2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n507), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n455), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n453), .A2(new_n448), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT35), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n586), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n575), .A2(new_n576), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n369), .B1(new_n614), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT11), .B(G169gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(G113gat), .B(G141gat), .Z(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n234), .A2(new_n235), .ZN(new_n631));
  AOI211_X1 g430(.A(KEYINPUT17), .B(new_n219), .C1(new_n233), .C2(new_n227), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n301), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n234), .B2(new_n301), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT97), .B(new_n301), .C1(new_n631), .C2(new_n632), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n635), .A2(KEYINPUT18), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n639));
  INV_X1    g438(.A(new_n301), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n230), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n234), .A2(new_n301), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n636), .B(KEYINPUT13), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n231), .B2(new_n236), .ZN(new_n647));
  INV_X1    g446(.A(new_n634), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n637), .B(new_n636), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n639), .B1(new_n638), .B2(new_n645), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n630), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n651), .A2(new_n629), .A3(new_n645), .A4(new_n638), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n624), .A2(KEYINPUT110), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT110), .B1(new_n624), .B2(new_n659), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n610), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(new_n662), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n621), .B1(new_n668), .B2(new_n660), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT111), .B1(new_n669), .B2(new_n300), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT111), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(G8gat), .C1(new_n663), .C2(new_n621), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NOR2_X1   g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n621), .B(new_n675), .C1(new_n668), .C2(new_n660), .ZN(new_n676));
  NAND2_X1  g475(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n675), .ZN(new_n679));
  AND4_X1   g478(.A1(new_n674), .A2(new_n669), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n673), .B1(new_n678), .B2(new_n680), .ZN(G1325gat));
  AOI21_X1  g480(.A(G15gat), .B1(new_n664), .B2(new_n615), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n455), .A2(KEYINPUT112), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n451), .A2(new_n454), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n663), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n687), .B2(G15gat), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n663), .A2(new_n612), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  AOI21_X1  g490(.A(new_n272), .B1(new_n614), .B2(new_n623), .ZN(new_n692));
  INV_X1    g491(.A(new_n659), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n367), .A2(new_n693), .A3(new_n319), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(G29gat), .A3(new_n610), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n686), .B1(new_n603), .B2(new_n613), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n623), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n271), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n702), .B2(new_n692), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n694), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n610), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n695), .A2(G36gat), .A3(new_n621), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT46), .ZN(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n705), .B2(new_n621), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1329gat));
  NAND3_X1  g510(.A1(new_n704), .A2(G43gat), .A3(new_n694), .ZN(new_n712));
  INV_X1    g511(.A(new_n615), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n695), .A2(new_n713), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n712), .A2(new_n686), .B1(G43gat), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g515(.A(G50gat), .B1(new_n705), .B2(new_n612), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n612), .B1(new_n695), .B2(KEYINPUT115), .ZN(new_n719));
  INV_X1    g518(.A(G50gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n719), .B(new_n720), .C1(KEYINPUT115), .C2(new_n695), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n717), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  AOI21_X1  g523(.A(new_n659), .B1(new_n700), .B2(new_n623), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n321), .A2(new_n367), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n665), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n621), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n727), .B2(new_n686), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n727), .A2(G71gat), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n615), .B(KEYINPUT116), .Z(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g540(.A1(new_n728), .A2(new_n507), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n659), .A2(new_n319), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n704), .A2(new_n367), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n248), .A3(new_n610), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n272), .B1(new_n700), .B2(new_n623), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n747), .A2(new_n748), .A3(new_n744), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n744), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n665), .A3(new_n367), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n746), .B1(new_n248), .B2(new_n752), .ZN(G1336gat));
  NAND4_X1  g552(.A1(new_n704), .A2(new_n622), .A3(new_n367), .A4(new_n744), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  INV_X1    g554(.A(new_n750), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n748), .A3(new_n744), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(new_n249), .A3(new_n367), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n621), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n754), .A2(G92gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n761), .B(new_n762), .C1(new_n621), .C2(new_n758), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n745), .B2(new_n686), .ZN(new_n765));
  INV_X1    g564(.A(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n766), .A3(new_n367), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n713), .B2(new_n767), .ZN(G1338gat));
  NAND4_X1  g567(.A1(new_n704), .A2(new_n507), .A3(new_n367), .A4(new_n744), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(G106gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n751), .A2(new_n771), .A3(new_n507), .A4(new_n367), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  INV_X1    g575(.A(new_n319), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n345), .A2(new_n347), .A3(new_n341), .A4(new_n348), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n357), .A2(KEYINPUT107), .A3(new_n341), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n327), .B1(new_n361), .B2(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n778), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n780), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT54), .B(new_n787), .C1(new_n352), .C2(new_n358), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n786), .A2(new_n659), .A3(new_n359), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n658), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n655), .A2(new_n656), .ZN(new_n792));
  INV_X1    g591(.A(new_n628), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n643), .A2(new_n644), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n635), .A2(new_n637), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n636), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n359), .A2(KEYINPUT109), .A3(new_n362), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT109), .B1(new_n359), .B2(new_n362), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n271), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n789), .A2(new_n359), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n788), .B2(new_n784), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n793), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n657), .B2(new_n658), .ZN(new_n805));
  NOR4_X1   g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n272), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n777), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n321), .A2(new_n368), .A3(new_n693), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n622), .A2(new_n610), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n618), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n693), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n659), .A2(new_n416), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT119), .Z(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n814), .B2(new_n817), .ZN(G1340gat));
  INV_X1    g617(.A(new_n814), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n413), .A3(new_n367), .ZN(new_n820));
  OAI21_X1  g619(.A(G120gat), .B1(new_n814), .B2(new_n368), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n822), .B(new_n823), .ZN(G1341gat));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n319), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g625(.A1(new_n814), .A2(new_n272), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n828));
  XOR2_X1   g627(.A(KEYINPUT56), .B(G134gat), .Z(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(G1343gat));
  NOR3_X1   g629(.A1(new_n810), .A2(new_n811), .A3(new_n612), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n809), .ZN(new_n834));
  INV_X1    g633(.A(new_n806), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n659), .A2(new_n789), .A3(new_n359), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT121), .B1(new_n783), .B2(new_n785), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n788), .A2(new_n839), .A3(new_n784), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n778), .A3(new_n840), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n837), .A2(new_n841), .B1(new_n367), .B2(new_n797), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n835), .B1(new_n842), .B2(new_n271), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n834), .B1(new_n843), .B2(new_n777), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT57), .B1(new_n844), .B2(new_n612), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n813), .A2(new_n686), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n833), .A2(new_n845), .A3(new_n659), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  INV_X1    g648(.A(G141gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n850), .A3(new_n659), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n851), .B2(KEYINPUT122), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n849), .B(new_n851), .C1(KEYINPUT122), .C2(new_n853), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(G148gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n847), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT59), .B(new_n858), .C1(new_n859), .C2(new_n368), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n836), .A2(new_n803), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n805), .B1(new_n365), .B2(new_n366), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n272), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n319), .B1(new_n864), .B2(new_n835), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n865), .B2(new_n834), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(KEYINPUT57), .A3(new_n507), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n840), .A2(new_n778), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n839), .B1(new_n788), .B2(new_n784), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n800), .B1(new_n872), .B2(new_n836), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n806), .B1(new_n873), .B2(new_n272), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n809), .B1(new_n874), .B2(new_n319), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n507), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n868), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n812), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n507), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(KEYINPUT59), .A3(new_n367), .A4(new_n847), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n833), .A2(new_n847), .A3(new_n845), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n368), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(KEYINPUT59), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n861), .B1(new_n883), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g683(.A(new_n468), .B1(new_n859), .B2(new_n777), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n881), .A2(new_n777), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n468), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(new_n469), .B1(new_n859), .B2(new_n272), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n881), .A2(new_n272), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n469), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n810), .A2(new_n811), .A3(new_n665), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n621), .A2(new_n616), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT124), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n381), .A3(new_n659), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n739), .A2(new_n507), .A3(new_n621), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n693), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n896), .B2(new_n367), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n899), .A2(new_n323), .A3(new_n368), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1349gat));
  OAI21_X1  g703(.A(new_n389), .B1(new_n899), .B2(new_n777), .ZN(new_n905));
  INV_X1    g704(.A(new_n896), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n777), .A2(new_n401), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n377), .A3(new_n271), .A4(new_n895), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT125), .ZN(new_n911));
  OAI21_X1  g710(.A(G190gat), .B1(new_n899), .B2(new_n272), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT61), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n912), .A2(KEYINPUT61), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n686), .A2(new_n610), .A3(new_n622), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n877), .B2(new_n878), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G197gat), .B1(new_n919), .B2(new_n693), .ZN(new_n920));
  INV_X1    g719(.A(new_n917), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n866), .A2(new_n507), .A3(new_n921), .A4(new_n867), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  INV_X1    g722(.A(G197gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n659), .A4(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n920), .B1(new_n927), .B2(new_n928), .ZN(G1352gat));
  NOR3_X1   g728(.A1(new_n922), .A2(G204gat), .A3(new_n368), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n368), .B(new_n917), .C1(new_n877), .C2(new_n878), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n325), .ZN(G1353gat));
  NAND4_X1  g734(.A1(new_n923), .A2(new_n309), .A3(new_n319), .A4(new_n925), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n937), .B(new_n309), .C1(new_n918), .C2(new_n319), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n832), .B1(new_n844), .B2(new_n612), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n831), .A2(KEYINPUT57), .B1(new_n939), .B2(KEYINPUT123), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n868), .A2(new_n869), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n319), .B(new_n921), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n936), .B1(new_n938), .B2(new_n943), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n919), .B2(new_n272), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n925), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n271), .A2(new_n458), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1355gat));
endmodule


