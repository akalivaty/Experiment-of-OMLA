//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n221), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G97), .B(G107), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  INV_X1    g0051(.A(new_n216), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n250), .A2(G226), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT66), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n261), .B1(new_n262), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT10), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n268), .A2(new_n269), .B1(KEYINPUT69), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n258), .B2(new_n267), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n216), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n206), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G50), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G50), .B2(new_n276), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT64), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n207), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT64), .A2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G33), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n285), .A2(new_n289), .A3(G33), .A4(new_n286), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n283), .B1(new_n297), .B2(new_n279), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT9), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n274), .A2(new_n275), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n275), .B1(new_n274), .B2(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n268), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G179), .B2(new_n268), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n256), .A2(new_n247), .A3(G274), .ZN(new_n306));
  INV_X1    g0106(.A(G244), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n249), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n309));
  INV_X1    g0109(.A(G107), .ZN(new_n310));
  INV_X1    g0110(.A(G238), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n309), .B1(new_n310), .B2(new_n259), .C1(new_n263), .C2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n308), .B1(new_n312), .B2(new_n266), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G190), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n272), .B2(new_n313), .ZN(new_n315));
  INV_X1    g0115(.A(new_n279), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  NAND2_X1  g0117(.A1(new_n291), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n288), .A2(KEYINPUT68), .A3(new_n290), .A4(new_n317), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT64), .B(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n293), .A2(new_n295), .B1(new_n322), .B2(G77), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n316), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n281), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n262), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n280), .A2(new_n327), .B1(new_n262), .B2(new_n277), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n315), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(new_n329), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n313), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G169), .B2(new_n313), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n305), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  OAI211_X1 g0143(.A(G232), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(G226), .B(new_n260), .C1(new_n342), .C2(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT71), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G33), .A3(G97), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n266), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT72), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n306), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n256), .A2(new_n247), .A3(KEYINPUT72), .A4(G274), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n247), .A2(G238), .A3(new_n248), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT13), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n352), .A2(new_n357), .A3(new_n360), .A4(new_n354), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(KEYINPUT73), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n366), .A3(KEYINPUT13), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n365), .A2(new_n367), .A3(G179), .A4(new_n361), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n369), .A3(G169), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT12), .B1(new_n276), .B2(G68), .ZN(new_n372));
  OR3_X1    g0172(.A1(new_n276), .A2(KEYINPUT12), .A3(G68), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n326), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n372), .A2(new_n373), .B1(new_n280), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n288), .A2(G77), .A3(new_n290), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n374), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n279), .ZN(new_n381));
  INV_X1    g0181(.A(new_n377), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n316), .B(new_n382), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n376), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n272), .B1(new_n359), .B2(new_n361), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n384), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n358), .A2(new_n366), .A3(KEYINPUT13), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n366), .B1(new_n358), .B2(KEYINPUT13), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n361), .A2(G190), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND4_X1   g0194(.A1(new_n389), .A2(new_n365), .A3(new_n367), .A4(new_n393), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n292), .A2(new_n326), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n280), .B1(new_n277), .B2(new_n292), .ZN(new_n400));
  AND2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n295), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(KEYINPUT3), .A2(G33), .ZN(new_n406));
  NAND2_X1  g0206(.A1(KEYINPUT3), .A2(G33), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n207), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n322), .A2(new_n259), .A3(KEYINPUT7), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n405), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n279), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT7), .B1(new_n322), .B2(new_n259), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n342), .A2(new_n343), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n207), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(G68), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n420), .B2(new_n405), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n400), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(G223), .B(new_n260), .C1(new_n342), .C2(new_n343), .ZN(new_n423));
  OAI211_X1 g0223(.A(G226), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n266), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n250), .A2(G232), .B1(new_n253), .B2(new_n256), .ZN(new_n428));
  AOI21_X1  g0228(.A(G200), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n269), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n398), .B1(new_n422), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n400), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n420), .A2(new_n405), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n414), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n374), .B1(new_n408), .B2(KEYINPUT7), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n215), .A2(new_n417), .A3(new_n418), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n404), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n316), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n427), .A2(new_n428), .A3(G179), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n302), .B1(new_n427), .B2(new_n428), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT18), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n427), .A2(new_n428), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G169), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n332), .B2(new_n445), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n422), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n427), .A2(new_n428), .A3(new_n269), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n430), .B2(G200), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n432), .A2(new_n444), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n397), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n341), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n255), .A2(G1), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(G274), .A3(new_n247), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n266), .B1(new_n457), .B2(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(KEYINPUT82), .A3(G270), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G270), .A3(new_n247), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n459), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n259), .A2(new_n471), .A3(G264), .A4(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n417), .A2(G303), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n259), .A2(G257), .A3(new_n260), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n475), .A2(new_n476), .A3(new_n266), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n475), .B2(new_n266), .ZN(new_n478));
  OAI211_X1 g0278(.A(G190), .B(new_n468), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n277), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n276), .A2(new_n482), .A3(new_n216), .A4(new_n278), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n215), .B(new_n485), .C1(G33), .C2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n278), .A2(new_n216), .B1(G20), .B2(new_n480), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT82), .B1(new_n460), .B2(G270), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n465), .A2(new_n466), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n458), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n475), .A2(new_n266), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n475), .A2(new_n476), .A3(new_n266), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n479), .B(new_n493), .C1(new_n500), .C2(new_n272), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n491), .A2(new_n492), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(G169), .C1(new_n503), .C2(new_n484), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT21), .B1(new_n493), .B2(new_n302), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT21), .B1(new_n493), .B2(new_n332), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n500), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n501), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n464), .A2(new_n247), .ZN(new_n511));
  INV_X1    g0311(.A(G257), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n458), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(new_n260), .C1(new_n342), .C2(new_n343), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n485), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n519), .B2(new_n266), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n332), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n266), .ZN(new_n522));
  INV_X1    g0322(.A(new_n513), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n302), .ZN(new_n525));
  NOR4_X1   g0325(.A1(new_n262), .A2(KEYINPUT78), .A3(G20), .A4(G33), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n295), .B2(G77), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n310), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  XNOR2_X1  g0330(.A(G97), .B(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n529), .B1(new_n533), .B2(new_n215), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n416), .A2(G107), .A3(new_n419), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(KEYINPUT79), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n416), .A2(new_n537), .A3(G107), .A4(new_n419), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n316), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n483), .A2(G97), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n276), .A2(new_n486), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n521), .B(new_n525), .C1(new_n539), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n522), .A2(new_n269), .A3(new_n523), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G200), .B2(new_n520), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n549));
  INV_X1    g0349(.A(new_n534), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n538), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n545), .B1(new_n551), .B2(new_n279), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n288), .A2(G97), .A3(new_n290), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n215), .ZN(new_n558));
  XNOR2_X1  g0358(.A(KEYINPUT81), .B(G87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n486), .A3(new_n310), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n417), .A2(new_n322), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n558), .A2(new_n560), .B1(new_n561), .B2(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n279), .ZN(new_n564));
  INV_X1    g0364(.A(new_n317), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n277), .ZN(new_n566));
  INV_X1    g0366(.A(new_n483), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n317), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n247), .A2(G274), .A3(new_n457), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n206), .A2(G45), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n247), .A2(G250), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G244), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n574));
  OAI211_X1 g0374(.A(G238), .B(new_n260), .C1(new_n342), .C2(new_n343), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G116), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n577), .B2(new_n266), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G179), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n302), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n269), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G200), .B2(new_n578), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n567), .A2(G87), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n564), .A3(new_n566), .A4(new_n584), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n546), .A2(new_n553), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n464), .A2(G264), .A3(new_n247), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G250), .A2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n512), .B2(G1698), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n259), .B1(G33), .B2(G294), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n266), .B1(new_n591), .B2(KEYINPUT86), .ZN(new_n592));
  OR2_X1    g0392(.A1(G250), .A2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n512), .A2(G1698), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(new_n342), .C2(new_n343), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n458), .B(new_n588), .C1(new_n592), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT88), .B1(new_n600), .B2(G190), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n272), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n247), .B1(new_n597), .B2(new_n598), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n587), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n269), .A4(new_n458), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n215), .A2(new_n259), .A3(G87), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT22), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT24), .ZN(new_n611));
  NAND2_X1  g0411(.A1(KEYINPUT23), .A2(G107), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(G20), .ZN(new_n614));
  OR2_X1    g0414(.A1(KEYINPUT23), .A2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n322), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n611), .B1(new_n610), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n279), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n277), .A2(new_n310), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT25), .ZN(new_n623));
  XOR2_X1   g0423(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n567), .B2(G107), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n600), .A2(G169), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n332), .C2(new_n600), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n600), .A2(new_n332), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n302), .B1(new_n605), .B2(new_n458), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT87), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n510), .A2(new_n586), .A3(new_n627), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n455), .A2(new_n636), .ZN(G372));
  AND2_X1   g0437(.A1(new_n581), .A2(new_n585), .ZN(new_n638));
  INV_X1    g0438(.A(new_n546), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(KEYINPUT90), .A3(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(KEYINPUT89), .A3(new_n646), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n643), .A2(new_n644), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n586), .A2(new_n627), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n507), .A2(new_n509), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n632), .A2(new_n633), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n628), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n652), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n581), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n455), .B1(new_n651), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n444), .A2(new_n449), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n387), .A2(new_n384), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n365), .A2(new_n393), .A3(new_n367), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT74), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n392), .A2(new_n389), .A3(new_n393), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n335), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n386), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n432), .A2(new_n452), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n662), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n300), .A2(new_n301), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n304), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n661), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n215), .A2(new_n206), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n653), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT91), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n628), .A2(new_n681), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n635), .A2(new_n627), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n635), .B2(new_n682), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n657), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n682), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n682), .A2(new_n493), .ZN(new_n692));
  MUX2_X1   g0492(.A(new_n510), .B(new_n653), .S(new_n692), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n687), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n210), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n206), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n560), .A2(G116), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n700), .A2(new_n701), .B1(new_n220), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT93), .B1(new_n654), .B2(new_n635), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n652), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n654), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n659), .B1(new_n641), .B2(new_n647), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n681), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n681), .B1(new_n651), .B2(new_n660), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n710), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n636), .A2(KEYINPUT31), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n332), .B(new_n573), .C1(new_n266), .C2(new_n577), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n520), .A3(new_n605), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n505), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT92), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT92), .B(new_n715), .C1(new_n505), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n505), .A2(new_n717), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n578), .A2(G179), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n600), .A2(new_n524), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n724), .A2(KEYINPUT30), .B1(new_n505), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n681), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n714), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n727), .A2(new_n718), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n681), .A2(KEYINPUT31), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n711), .A2(new_n713), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n703), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n322), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n700), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n695), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n693), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n698), .A2(new_n417), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G355), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G116), .B2(new_n210), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n698), .A2(new_n259), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n255), .B2(new_n220), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n241), .A2(new_n255), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT94), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n755), .B2(G20), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(KEYINPUT94), .A3(new_n207), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n216), .B1(G20), .B2(new_n302), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n742), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n215), .A2(new_n332), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n269), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G50), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n272), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n322), .A2(new_n269), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G107), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n767), .A2(G20), .A3(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n559), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n417), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n766), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n269), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n763), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n778), .A2(G77), .B1(new_n781), .B2(G58), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n322), .A2(new_n269), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n215), .B1(new_n332), .B2(new_n779), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n782), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n764), .A2(G190), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n775), .B(new_n791), .C1(G68), .C2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n792), .A2(new_n796), .B1(new_n781), .B2(G322), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n777), .A2(new_n799), .B1(new_n800), .B2(new_n768), .ZN(new_n801));
  INV_X1    g0601(.A(new_n784), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G329), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n417), .B1(new_n804), .B2(new_n771), .C1(new_n788), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G326), .B2(new_n765), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n798), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n794), .A2(new_n795), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n762), .B1(new_n809), .B2(new_n759), .ZN(new_n810));
  INV_X1    g0610(.A(new_n758), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n693), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n331), .A2(new_n682), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n668), .B1(new_n330), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n335), .A2(new_n682), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n712), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n742), .B1(new_n819), .B2(new_n734), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n734), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n759), .A2(new_n754), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n741), .B1(new_n262), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n789), .A2(G58), .B1(new_n802), .B2(G132), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n769), .A2(G68), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n417), .B1(new_n772), .B2(G50), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n778), .A2(G159), .B1(new_n781), .B2(G143), .ZN(new_n828));
  INV_X1    g0628(.A(new_n792), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(new_n765), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n827), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n790), .B1(new_n780), .B2(new_n805), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT97), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n800), .A2(new_n829), .B1(new_n832), .B2(new_n804), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n417), .B1(new_n310), .B2(new_n771), .C1(new_n784), .C2(new_n799), .ZN(new_n840));
  INV_X1    g0640(.A(G87), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n777), .A2(new_n480), .B1(new_n841), .B2(new_n768), .ZN(new_n842));
  OR3_X1    g0642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n836), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n759), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(KEYINPUT98), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n823), .B1(new_n755), .B2(new_n818), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n821), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n739), .A2(new_n206), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n455), .B1(new_n711), .B2(new_n713), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n674), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  INV_X1    g0654(.A(new_n817), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n712), .B2(new_n818), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n405), .B1(new_n410), .B2(new_n411), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n414), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n433), .B1(new_n859), .B2(new_n439), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT100), .B1(new_n860), .B2(new_n679), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n438), .A2(new_n415), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n400), .B1(new_n413), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT100), .ZN(new_n864));
  INV_X1    g0664(.A(new_n679), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n440), .A2(new_n451), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n443), .B2(new_n860), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n422), .A2(new_n447), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n422), .A2(new_n865), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n868), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n453), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT101), .B1(new_n453), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n875), .B(KEYINPUT38), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n385), .A2(new_n681), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n386), .A2(new_n396), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n386), .B2(new_n396), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n857), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n453), .A2(new_n867), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n453), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n893), .B2(new_n875), .ZN(new_n894));
  INV_X1    g0694(.A(new_n881), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT39), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n386), .A2(new_n681), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n871), .A2(new_n872), .A3(new_n868), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n440), .A2(new_n679), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n900), .A2(new_n874), .B1(new_n453), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n881), .B1(KEYINPUT38), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n897), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n662), .A2(new_n679), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n888), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n854), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(G330), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n716), .A2(new_n520), .A3(new_n605), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n500), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT92), .B1(new_n912), .B2(new_n715), .ZN(new_n913));
  INV_X1    g0713(.A(new_n721), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n727), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n732), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n455), .B1(new_n730), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n816), .A2(new_n817), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n385), .B(new_n681), .C1(new_n667), .C2(new_n371), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n386), .A2(new_n396), .A3(new_n883), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n918), .B(new_n732), .C1(new_n722), .C2(new_n727), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT103), .B1(new_n915), .B2(new_n916), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n636), .A2(KEYINPUT31), .B1(new_n681), .B2(new_n728), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n896), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n730), .A2(new_n921), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n882), .A2(new_n936), .A3(new_n927), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n818), .B1(new_n884), .B2(new_n885), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n730), .B2(new_n921), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n935), .A2(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n910), .B1(new_n922), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n922), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n851), .B1(new_n909), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n909), .B2(new_n945), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n219), .A2(new_n262), .A3(new_n401), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n374), .A2(G50), .ZN(new_n949));
  OAI211_X1 g0749(.A(G1), .B(new_n738), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n533), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n217), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n950), .A3(new_n956), .ZN(G367));
  OAI211_X1 g0757(.A(new_n546), .B(new_n553), .C1(new_n552), .C2(new_n682), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n546), .B2(new_n682), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n689), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT42), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(KEYINPUT106), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n546), .B1(new_n962), .B2(new_n635), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n961), .B1(new_n682), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n564), .A2(new_n566), .A3(new_n584), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n681), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n638), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT105), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT105), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n967), .A2(new_n581), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n964), .A2(new_n965), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT107), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n972), .B(KEYINPUT43), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n964), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n696), .A2(new_n962), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n740), .A2(G1), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n691), .A2(new_n959), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT45), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n691), .A2(new_n959), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n696), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n694), .B(new_n687), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n684), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n735), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n736), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n699), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n982), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n981), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n973), .A2(new_n758), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n749), .A2(new_n237), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n760), .B1(new_n210), .B2(new_n565), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n742), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n832), .A2(new_n799), .B1(new_n804), .B2(new_n780), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n788), .A2(new_n310), .B1(new_n486), .B2(new_n768), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n777), .A2(new_n800), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G317), .C2(new_n802), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n772), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n771), .B2(new_n480), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n417), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G294), .B2(new_n792), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n788), .A2(new_n374), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n202), .A2(new_n777), .B1(new_n780), .B2(new_n830), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G137), .C2(new_n802), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n768), .A2(new_n262), .ZN(new_n1018));
  INV_X1    g0818(.A(G58), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n259), .B1(new_n771), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n765), .C2(G143), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(new_n1021), .C1(new_n785), .C2(new_n829), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1002), .B1(new_n1024), .B2(new_n759), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n999), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n998), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n990), .A2(new_n982), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT109), .Z(new_n1031));
  NOR2_X1   g0831(.A1(new_n687), .A2(new_n811), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n234), .A2(new_n255), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n701), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1033), .A2(new_n748), .B1(new_n1034), .B2(new_n745), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n255), .B1(new_n374), .B2(new_n262), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n293), .B2(new_n202), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n292), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1035), .A2(new_n1040), .B1(G107), .B2(new_n210), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n741), .B1(new_n1041), .B2(new_n760), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT110), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n759), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n778), .A2(G303), .B1(new_n781), .B2(G317), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n765), .A2(G322), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n799), .C2(new_n829), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n789), .A2(G283), .B1(new_n772), .B2(G294), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n768), .A2(new_n480), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n259), .B(new_n1056), .C1(G326), .C2(new_n802), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n788), .A2(new_n565), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n777), .A2(new_n374), .B1(new_n830), .B2(new_n784), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G50), .C2(new_n781), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n259), .B1(new_n262), .B2(new_n771), .C1(new_n768), .C2(new_n486), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n293), .B2(new_n792), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n785), .C2(new_n832), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1044), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1043), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT111), .B1(new_n991), .B2(new_n735), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n991), .A2(KEYINPUT111), .A3(new_n735), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n699), .C1(new_n735), .C2(new_n991), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1031), .B1(new_n1032), .B2(new_n1066), .C1(new_n1067), .C2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n699), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n988), .B2(new_n992), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n992), .B2(new_n988), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n749), .A2(new_n244), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n760), .B1(new_n486), .B2(new_n210), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n742), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT112), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n765), .A2(G317), .B1(new_n781), .B2(G311), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  OAI211_X1 g0879(.A(new_n770), .B(new_n417), .C1(new_n800), .C2(new_n771), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n789), .A2(G116), .B1(new_n802), .B2(G322), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n805), .B2(new_n777), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(G303), .C2(new_n792), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n765), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  OAI221_X1 g0885(.A(new_n259), .B1(new_n374), .B2(new_n771), .C1(new_n768), .C2(new_n841), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n802), .A2(G143), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n262), .B2(new_n788), .C1(new_n292), .C2(new_n777), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G50), .C2(new_n792), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1079), .A2(new_n1083), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1077), .B1(new_n1090), .B2(new_n1044), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n962), .B2(new_n758), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n988), .B2(new_n982), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1073), .A2(new_n1093), .ZN(G390));
  INV_X1    g0894(.A(new_n898), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n856), .B2(new_n886), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n897), .A2(new_n905), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n709), .A2(new_n816), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n887), .B1(new_n1098), .B2(new_n855), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n903), .A2(new_n1095), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1096), .A2(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n733), .A2(G330), .A3(new_n818), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(new_n886), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n936), .A2(G330), .A3(new_n927), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G1), .B2(new_n740), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1097), .A2(new_n754), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n772), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n778), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n789), .A2(G159), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n202), .A2(new_n768), .B1(new_n784), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n417), .B(new_n1116), .C1(G132), .C2(new_n781), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G128), .A2(new_n765), .B1(new_n792), .B2(G137), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n825), .B(new_n417), .C1(new_n841), .C2(new_n771), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G107), .B2(new_n792), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n778), .A2(G97), .B1(new_n789), .B2(G77), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n781), .A2(G116), .B1(G294), .B2(new_n802), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n765), .A2(G283), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1044), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n741), .B(new_n1126), .C1(new_n292), .C2(new_n822), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1107), .B1(new_n1108), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n936), .A2(G330), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n455), .A2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n852), .A2(new_n1130), .A3(new_n674), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1098), .A2(new_n855), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n886), .B1(new_n1129), .B2(new_n924), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1103), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1129), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1102), .A2(new_n886), .B1(new_n927), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n856), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1071), .B1(new_n1106), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1106), .B2(new_n1138), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1128), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(new_n908), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n298), .A2(new_n679), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT55), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n305), .B(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(G330), .B1(new_n941), .B2(new_n932), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n934), .B(KEYINPUT40), .C1(new_n940), .C2(new_n882), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT104), .B1(new_n937), .B2(new_n923), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT115), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n935), .A2(new_n938), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT115), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n1150), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(KEYINPUT115), .B(new_n1149), .C1(new_n935), .C2(new_n938), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1147), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1142), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT116), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1156), .B1(new_n1155), .B2(new_n1150), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1147), .B1(new_n1163), .B2(new_n1159), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1148), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n908), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1162), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(KEYINPUT116), .A3(new_n1142), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1131), .B1(new_n1106), .B2(new_n1138), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT119), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT117), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1166), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1164), .A2(KEYINPUT117), .A3(new_n908), .A4(new_n1165), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT118), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1168), .B2(new_n1142), .ZN(new_n1179));
  AOI211_X1 g0979(.A(KEYINPUT118), .B(new_n908), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1176), .B(new_n1177), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1170), .A2(KEYINPUT57), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1071), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1171), .A2(new_n1184), .A3(new_n1172), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1174), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1167), .A2(new_n982), .A3(new_n1169), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n741), .B1(new_n202), .B2(new_n822), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n417), .A2(new_n254), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n772), .B2(G77), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n1019), .B2(new_n768), .C1(new_n800), .C2(new_n784), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT113), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n781), .A2(G107), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1015), .B1(new_n317), .B2(new_n778), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G97), .A2(new_n792), .B1(new_n765), .B2(G116), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n781), .A2(G128), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n778), .A2(G137), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n830), .B2(new_n788), .C1(new_n771), .C2(new_n1111), .ZN(new_n1202));
  INV_X1    g1002(.A(G132), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1115), .A2(new_n832), .B1(new_n829), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n769), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1189), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n1198), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1188), .B1(new_n1044), .B2(new_n1214), .C1(new_n1147), .C2(new_n755), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1187), .A2(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1186), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(G375));
  OR2_X1    g1018(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n996), .A3(new_n1138), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1137), .A2(new_n982), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n741), .B1(new_n374), .B2(new_n822), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT120), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n777), .A2(new_n830), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n780), .A2(new_n831), .B1(new_n788), .B2(new_n202), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(G128), .C2(new_n802), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n259), .B1(new_n785), .B2(new_n771), .C1(new_n768), .C2(new_n1019), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n792), .B2(new_n1112), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n1203), .C2(new_n832), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1059), .B1(G283), .B2(new_n781), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G116), .A2(new_n792), .B1(new_n765), .B2(G294), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n259), .B(new_n1018), .C1(G97), .C2(new_n772), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n778), .A2(G107), .B1(G303), .B2(new_n802), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1223), .B1(new_n1236), .B2(new_n759), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n887), .B2(new_n755), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1221), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1220), .A2(new_n1239), .ZN(G381));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n849), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1242), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1028), .A3(new_n1244), .A4(new_n1217), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(G407));
  NAND3_X1  g1046(.A1(new_n1217), .A2(new_n680), .A3(new_n1244), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G407), .A2(G213), .A3(new_n1247), .ZN(G409));
  XNOR2_X1  g1048(.A(G393), .B(new_n813), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1028), .A2(G390), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1241), .B1(new_n998), .B2(new_n1027), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1250), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI211_X1 g1055(.A(KEYINPUT124), .B(new_n1249), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1239), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1219), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(new_n1071), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1219), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1258), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(G384), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n680), .A2(G213), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G2897), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1264), .B(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1186), .A2(G378), .A3(new_n1216), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT123), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1186), .A2(KEYINPUT123), .A3(G378), .A4(new_n1216), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1181), .A2(new_n982), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n1215), .C1(new_n995), .C2(new_n1171), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1270), .A2(new_n1271), .B1(new_n1244), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1274), .B2(new_n1265), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1244), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1265), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1264), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1277), .A2(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1274), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1278), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1257), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1282), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1276), .A3(new_n1275), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1257), .B1(new_n1285), .B2(KEYINPUT63), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1257), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1286), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1276), .B(new_n1275), .C1(new_n1285), .C2(new_n1278), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1293), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(G405));
  NOR2_X1   g1100(.A1(new_n1217), .A2(G378), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT126), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1279), .ZN(new_n1303));
  OR3_X1    g1103(.A1(new_n1302), .A2(new_n1282), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1282), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1294), .ZN(G402));
endmodule


