

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767;

  XNOR2_X1 U375 ( .A(G104), .B(G143), .ZN(n413) );
  XNOR2_X2 U376 ( .A(n436), .B(n435), .ZN(n473) );
  XNOR2_X2 U377 ( .A(n602), .B(n601), .ZN(n686) );
  XOR2_X1 U378 ( .A(G137), .B(KEYINPUT4), .Z(n480) );
  XNOR2_X1 U379 ( .A(G128), .B(G137), .ZN(n493) );
  INV_X1 U380 ( .A(G953), .ZN(n449) );
  BUF_X1 U381 ( .A(G146), .Z(n368) );
  AND2_X2 U382 ( .A1(n421), .A2(n420), .ZN(n355) );
  NOR2_X2 U383 ( .A1(n759), .A2(n746), .ZN(n614) );
  XNOR2_X2 U384 ( .A(n403), .B(n394), .ZN(n759) );
  NOR2_X2 U385 ( .A1(n613), .A2(n736), .ZN(n598) );
  XNOR2_X2 U386 ( .A(n388), .B(n597), .ZN(n736) );
  XNOR2_X1 U387 ( .A(n573), .B(n444), .ZN(n553) );
  NAND2_X1 U388 ( .A1(n544), .A2(n516), .ZN(n747) );
  NOR2_X1 U389 ( .A1(n660), .A2(n473), .ZN(n397) );
  INV_X1 U390 ( .A(n368), .ZN(n390) );
  XNOR2_X1 U391 ( .A(n376), .B(n453), .ZN(n529) );
  NAND2_X1 U392 ( .A1(n553), .A2(n452), .ZN(n376) );
  XNOR2_X1 U393 ( .A(n397), .B(n439), .ZN(n526) );
  NOR2_X1 U394 ( .A1(n640), .A2(G902), .ZN(n385) );
  XNOR2_X1 U395 ( .A(n580), .B(n390), .ZN(n509) );
  XNOR2_X1 U396 ( .A(n482), .B(n391), .ZN(n580) );
  XNOR2_X1 U397 ( .A(n414), .B(G131), .ZN(n481) );
  XNOR2_X1 U398 ( .A(n456), .B(G134), .ZN(n482) );
  INV_X1 U399 ( .A(KEYINPUT72), .ZN(n414) );
  INV_X1 U400 ( .A(G125), .ZN(n426) );
  INV_X1 U401 ( .A(KEYINPUT86), .ZN(n371) );
  INV_X1 U402 ( .A(G478), .ZN(n384) );
  INV_X1 U403 ( .A(G902), .ZN(n489) );
  AND2_X1 U404 ( .A1(n373), .A2(n370), .ZN(n407) );
  XNOR2_X1 U405 ( .A(n372), .B(n371), .ZN(n370) );
  NAND2_X1 U406 ( .A1(n556), .A2(n555), .ZN(n372) );
  XNOR2_X1 U407 ( .A(n381), .B(KEYINPUT36), .ZN(n380) );
  NAND2_X1 U408 ( .A1(n365), .A2(n364), .ZN(n381) );
  INV_X1 U409 ( .A(n575), .ZN(n365) );
  XNOR2_X1 U410 ( .A(n523), .B(KEYINPUT112), .ZN(n575) );
  NAND2_X1 U411 ( .A1(n529), .A2(n477), .ZN(n367) );
  NOR2_X1 U412 ( .A1(n377), .A2(n596), .ZN(n589) );
  NOR2_X1 U413 ( .A1(n539), .A2(n538), .ZN(n542) );
  AND2_X1 U414 ( .A1(n532), .A2(n705), .ZN(n714) );
  BUF_X1 U415 ( .A(n572), .Z(n705) );
  XNOR2_X1 U416 ( .A(n572), .B(KEYINPUT93), .ZN(n377) );
  NOR2_X1 U417 ( .A1(n549), .A2(n382), .ZN(n522) );
  XNOR2_X1 U418 ( .A(n561), .B(n560), .ZN(n726) );
  INV_X1 U419 ( .A(n574), .ZN(n364) );
  AND2_X1 U420 ( .A1(n747), .A2(n749), .ZN(n723) );
  NAND2_X1 U421 ( .A1(n526), .A2(n724), .ZN(n573) );
  AND2_X1 U422 ( .A1(n516), .A2(n707), .ZN(n383) );
  XNOR2_X1 U423 ( .A(n711), .B(KEYINPUT6), .ZN(n596) );
  BUF_X1 U424 ( .A(n711), .Z(n366) );
  INV_X1 U425 ( .A(n534), .ZN(n544) );
  XNOR2_X1 U426 ( .A(n385), .B(n384), .ZN(n534) );
  XNOR2_X1 U427 ( .A(n408), .B(n472), .ZN(n543) );
  XNOR2_X1 U428 ( .A(n507), .B(n379), .ZN(n378) );
  XNOR2_X1 U429 ( .A(n509), .B(n488), .ZN(n653) );
  XNOR2_X1 U430 ( .A(n457), .B(n386), .ZN(n640) );
  OR2_X1 U431 ( .A1(n492), .A2(n646), .ZN(n457) );
  XNOR2_X1 U432 ( .A(n506), .B(n508), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n482), .B(n461), .ZN(n386) );
  XNOR2_X1 U434 ( .A(n438), .B(KEYINPUT96), .ZN(n439) );
  XNOR2_X1 U435 ( .A(n480), .B(n481), .ZN(n391) );
  XNOR2_X1 U436 ( .A(n692), .B(KEYINPUT75), .ZN(n507) );
  XNOR2_X1 U437 ( .A(n427), .B(G107), .ZN(n692) );
  XNOR2_X2 U438 ( .A(G119), .B(G110), .ZN(n494) );
  XNOR2_X1 U439 ( .A(G902), .B(KEYINPUT94), .ZN(n436) );
  XNOR2_X2 U440 ( .A(G104), .B(G110), .ZN(n427) );
  XNOR2_X1 U441 ( .A(n357), .B(n356), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n359), .B(n456), .ZN(n356) );
  XNOR2_X1 U443 ( .A(n358), .B(n360), .ZN(n357) );
  NAND2_X1 U444 ( .A1(n642), .A2(G224), .ZN(n358) );
  XNOR2_X1 U445 ( .A(n361), .B(G125), .ZN(n359) );
  XNOR2_X1 U446 ( .A(n362), .B(n363), .ZN(n360) );
  XNOR2_X2 U447 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n361) );
  XNOR2_X2 U448 ( .A(KEYINPUT83), .B(G146), .ZN(n362) );
  XNOR2_X2 U449 ( .A(KEYINPUT18), .B(KEYINPUT95), .ZN(n363) );
  XNOR2_X2 U450 ( .A(n428), .B(G953), .ZN(n642) );
  NOR2_X2 U451 ( .A1(n355), .A2(n632), .ZN(n417) );
  XNOR2_X2 U452 ( .A(n367), .B(n478), .ZN(n592) );
  BUF_X2 U453 ( .A(n642), .Z(n369) );
  NOR2_X1 U454 ( .A1(n559), .A2(n762), .ZN(n373) );
  XNOR2_X2 U455 ( .A(n374), .B(n392), .ZN(n579) );
  XNOR2_X2 U456 ( .A(n375), .B(KEYINPUT71), .ZN(n374) );
  XNOR2_X2 U457 ( .A(KEYINPUT10), .B(G140), .ZN(n375) );
  NOR2_X1 U458 ( .A1(n380), .A2(n377), .ZN(n762) );
  XNOR2_X1 U459 ( .A(n509), .B(n378), .ZN(n680) );
  NAND2_X1 U460 ( .A1(n544), .A2(n383), .ZN(n382) );
  INV_X1 U461 ( .A(n747), .ZN(n758) );
  XNOR2_X1 U462 ( .A(n387), .B(n507), .ZN(n434) );
  NAND2_X1 U463 ( .A1(n705), .A2(n389), .ZN(n388) );
  AND2_X1 U464 ( .A1(n596), .A2(n704), .ZN(n389) );
  XNOR2_X2 U465 ( .A(n426), .B(n368), .ZN(n392) );
  BUF_X1 U466 ( .A(n635), .Z(n393) );
  BUF_X1 U467 ( .A(n529), .Z(n530) );
  NOR2_X1 U468 ( .A1(n615), .A2(n723), .ZN(n617) );
  INV_X1 U469 ( .A(KEYINPUT15), .ZN(n435) );
  NOR2_X1 U470 ( .A1(G953), .A2(G237), .ZN(n483) );
  XNOR2_X1 U471 ( .A(G101), .B(KEYINPUT3), .ZN(n430) );
  XNOR2_X1 U472 ( .A(n469), .B(n409), .ZN(n671) );
  XNOR2_X1 U473 ( .A(n579), .B(n468), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n410) );
  INV_X1 U475 ( .A(KEYINPUT87), .ZN(n411) );
  NOR2_X1 U476 ( .A1(n620), .A2(n619), .ZN(n626) );
  XOR2_X1 U477 ( .A(KEYINPUT100), .B(KEYINPUT20), .Z(n474) );
  XOR2_X1 U478 ( .A(KEYINPUT12), .B(KEYINPUT105), .Z(n463) );
  XNOR2_X1 U479 ( .A(G113), .B(G122), .ZN(n462) );
  XNOR2_X1 U480 ( .A(n481), .B(n413), .ZN(n464) );
  NAND2_X1 U481 ( .A1(G234), .A2(G237), .ZN(n445) );
  XOR2_X1 U482 ( .A(KEYINPUT98), .B(KEYINPUT14), .Z(n446) );
  INV_X1 U483 ( .A(n530), .ZN(n613) );
  BUF_X1 U484 ( .A(n631), .Z(n636) );
  XNOR2_X1 U485 ( .A(KEYINPUT16), .B(G122), .ZN(n432) );
  XNOR2_X1 U486 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n454) );
  XNOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n495) );
  XNOR2_X1 U488 ( .A(G116), .B(G107), .ZN(n458) );
  NAND2_X1 U489 ( .A1(n671), .A2(n489), .ZN(n408) );
  XOR2_X1 U490 ( .A(G140), .B(G101), .Z(n508) );
  INV_X1 U491 ( .A(KEYINPUT42), .ZN(n396) );
  XNOR2_X1 U492 ( .A(n566), .B(n565), .ZN(n766) );
  NAND2_X1 U493 ( .A1(n530), .A2(n714), .ZN(n403) );
  XOR2_X1 U494 ( .A(n533), .B(KEYINPUT102), .Z(n394) );
  XNOR2_X1 U495 ( .A(KEYINPUT48), .B(KEYINPUT73), .ZN(n395) );
  XNOR2_X1 U496 ( .A(n396), .B(n571), .ZN(n767) );
  XNOR2_X1 U497 ( .A(n499), .B(n498), .ZN(n648) );
  NAND2_X2 U498 ( .A1(n700), .A2(KEYINPUT2), .ZN(n702) );
  NOR2_X2 U499 ( .A1(n635), .A2(n637), .ZN(n700) );
  AND2_X2 U500 ( .A1(n404), .A2(n425), .ZN(n631) );
  XNOR2_X1 U501 ( .A(n405), .B(n395), .ZN(n404) );
  NAND2_X1 U502 ( .A1(n416), .A2(KEYINPUT65), .ZN(n399) );
  NAND2_X1 U503 ( .A1(n398), .A2(n633), .ZN(n400) );
  NAND2_X1 U504 ( .A1(n399), .A2(n400), .ZN(n415) );
  INV_X1 U505 ( .A(n416), .ZN(n398) );
  NAND2_X1 U506 ( .A1(n419), .A2(n417), .ZN(n416) );
  BUF_X1 U507 ( .A(n594), .Z(n401) );
  XNOR2_X1 U508 ( .A(n423), .B(KEYINPUT32), .ZN(n594) );
  XNOR2_X1 U509 ( .A(n418), .B(KEYINPUT46), .ZN(n406) );
  OR2_X2 U510 ( .A1(n648), .A2(G902), .ZN(n505) );
  XNOR2_X1 U511 ( .A(n497), .B(n579), .ZN(n498) );
  NAND2_X1 U512 ( .A1(n402), .A2(n594), .ZN(n595) );
  XNOR2_X1 U513 ( .A(n402), .B(G110), .ZN(G12) );
  XNOR2_X2 U514 ( .A(n422), .B(KEYINPUT110), .ZN(n402) );
  NAND2_X1 U515 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U516 ( .A1(n603), .A2(n686), .ZN(n606) );
  NOR2_X1 U517 ( .A1(n608), .A2(n607), .ZN(n628) );
  NAND2_X1 U518 ( .A1(n756), .A2(n410), .ZN(n546) );
  NAND2_X1 U519 ( .A1(n723), .A2(KEYINPUT47), .ZN(n412) );
  NAND2_X2 U520 ( .A1(n415), .A2(n702), .ZN(n678) );
  NOR2_X2 U521 ( .A1(n766), .A2(n767), .ZN(n418) );
  INV_X1 U522 ( .A(n588), .ZN(n708) );
  XNOR2_X1 U523 ( .A(n611), .B(KEYINPUT113), .ZN(n539) );
  AND2_X2 U524 ( .A1(n704), .A2(n537), .ZN(n611) );
  NOR2_X2 U525 ( .A1(n588), .A2(n517), .ZN(n704) );
  NAND2_X1 U526 ( .A1(n634), .A2(n420), .ZN(n419) );
  XNOR2_X1 U527 ( .A(n629), .B(KEYINPUT45), .ZN(n634) );
  INV_X1 U528 ( .A(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U529 ( .A(n631), .B(n630), .ZN(n421) );
  NAND2_X1 U530 ( .A1(n592), .A2(n593), .ZN(n422) );
  NAND2_X1 U531 ( .A1(n592), .A2(n424), .ZN(n423) );
  AND2_X1 U532 ( .A1(n589), .A2(n588), .ZN(n424) );
  AND2_X1 U533 ( .A1(n765), .A2(n578), .ZN(n425) );
  AND2_X1 U534 ( .A1(n622), .A2(KEYINPUT76), .ZN(n623) );
  INV_X1 U535 ( .A(KEYINPUT80), .ZN(n630) );
  XNOR2_X1 U536 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U537 ( .A(KEYINPUT65), .ZN(n633) );
  BUF_X1 U538 ( .A(n660), .Z(n663) );
  INV_X1 U539 ( .A(KEYINPUT40), .ZN(n565) );
  XNOR2_X2 U540 ( .A(G128), .B(G143), .ZN(n456) );
  INV_X2 U541 ( .A(KEYINPUT64), .ZN(n428) );
  XNOR2_X2 U542 ( .A(G116), .B(G113), .ZN(n429) );
  XNOR2_X1 U543 ( .A(n429), .B(G119), .ZN(n431) );
  XNOR2_X1 U544 ( .A(n431), .B(n430), .ZN(n487) );
  INV_X1 U545 ( .A(n487), .ZN(n433) );
  XNOR2_X1 U546 ( .A(n433), .B(n432), .ZN(n693) );
  XNOR2_X1 U547 ( .A(n434), .B(n693), .ZN(n660) );
  INV_X1 U548 ( .A(G237), .ZN(n437) );
  NAND2_X1 U549 ( .A1(n437), .A2(n489), .ZN(n440) );
  NAND2_X1 U550 ( .A1(n440), .A2(G210), .ZN(n438) );
  NAND2_X1 U551 ( .A1(n440), .A2(G214), .ZN(n442) );
  INV_X1 U552 ( .A(KEYINPUT97), .ZN(n441) );
  XNOR2_X1 U553 ( .A(n442), .B(n441), .ZN(n724) );
  XNOR2_X1 U554 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n443), .B(KEYINPUT69), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U557 ( .A(KEYINPUT78), .B(n447), .Z(n448) );
  NAND2_X1 U558 ( .A1(G952), .A2(n448), .ZN(n734) );
  NOR2_X1 U559 ( .A1(n734), .A2(G953), .ZN(n521) );
  AND2_X1 U560 ( .A1(G902), .A2(n448), .ZN(n519) );
  NOR2_X1 U561 ( .A1(G898), .A2(n449), .ZN(n694) );
  NAND2_X1 U562 ( .A1(n519), .A2(n694), .ZN(n450) );
  XNOR2_X1 U563 ( .A(KEYINPUT99), .B(n450), .ZN(n451) );
  OR2_X1 U564 ( .A1(n521), .A2(n451), .ZN(n452) );
  INV_X1 U565 ( .A(KEYINPUT0), .ZN(n453) );
  NAND2_X1 U566 ( .A1(n642), .A2(G234), .ZN(n455) );
  XNOR2_X1 U567 ( .A(n455), .B(n454), .ZN(n492) );
  INV_X1 U568 ( .A(G217), .ZN(n646) );
  XNOR2_X1 U569 ( .A(n458), .B(KEYINPUT7), .ZN(n460) );
  XNOR2_X1 U570 ( .A(G122), .B(KEYINPUT9), .ZN(n459) );
  XNOR2_X1 U571 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U572 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U574 ( .A(KEYINPUT11), .B(KEYINPUT106), .Z(n467) );
  NAND2_X1 U575 ( .A1(G214), .A2(n483), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT13), .Z(n471) );
  XNOR2_X1 U578 ( .A(KEYINPUT107), .B(G475), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U580 ( .A1(n544), .A2(n543), .ZN(n721) );
  INV_X1 U581 ( .A(n473), .ZN(n632) );
  NAND2_X1 U582 ( .A1(n632), .A2(G234), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n475), .B(n474), .ZN(n500) );
  INV_X1 U584 ( .A(G221), .ZN(n491) );
  OR2_X1 U585 ( .A1(n500), .A2(n491), .ZN(n476) );
  XNOR2_X1 U586 ( .A(n476), .B(KEYINPUT21), .ZN(n517) );
  NOR2_X1 U587 ( .A1(n721), .A2(n517), .ZN(n477) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n478) );
  BUF_X1 U589 ( .A(n592), .Z(n479) );
  INV_X1 U590 ( .A(n479), .ZN(n515) );
  XOR2_X1 U591 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U592 ( .A1(n483), .A2(G210), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U594 ( .A1(n653), .A2(n489), .ZN(n490) );
  INV_X1 U595 ( .A(G472), .ZN(n651) );
  XNOR2_X2 U596 ( .A(n490), .B(n651), .ZN(n711) );
  OR2_X1 U597 ( .A1(n492), .A2(n491), .ZN(n499) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U600 ( .A(n500), .ZN(n501) );
  NAND2_X1 U601 ( .A1(n501), .A2(G217), .ZN(n503) );
  XNOR2_X1 U602 ( .A(KEYINPUT82), .B(KEYINPUT25), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X2 U604 ( .A(n505), .B(n504), .ZN(n588) );
  NOR2_X1 U605 ( .A1(n596), .A2(n588), .ZN(n513) );
  NAND2_X1 U606 ( .A1(n369), .A2(G227), .ZN(n506) );
  OR2_X1 U607 ( .A1(n680), .A2(G902), .ZN(n511) );
  XNOR2_X1 U608 ( .A(KEYINPUT74), .B(G469), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n511), .B(n510), .ZN(n537) );
  INV_X1 U610 ( .A(n537), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT68), .B(KEYINPUT1), .Z(n512) );
  XNOR2_X2 U612 ( .A(n551), .B(n512), .ZN(n572) );
  INV_X1 U613 ( .A(n572), .ZN(n590) );
  NAND2_X1 U614 ( .A1(n513), .A2(n590), .ZN(n514) );
  NOR2_X1 U615 ( .A1(n515), .A2(n514), .ZN(n616) );
  XOR2_X1 U616 ( .A(G101), .B(n616), .Z(G3) );
  INV_X1 U617 ( .A(n543), .ZN(n516) );
  INV_X1 U618 ( .A(n517), .ZN(n707) );
  NOR2_X1 U619 ( .A1(n369), .A2(G900), .ZN(n518) );
  AND2_X1 U620 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U621 ( .A1(n521), .A2(n520), .ZN(n538) );
  OR2_X1 U622 ( .A1(n708), .A2(n538), .ZN(n549) );
  NAND2_X1 U623 ( .A1(n596), .A2(n522), .ZN(n523) );
  NOR2_X1 U624 ( .A1(n575), .A2(n705), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n524), .A2(n724), .ZN(n525) );
  XNOR2_X1 U626 ( .A(KEYINPUT43), .B(n525), .ZN(n528) );
  BUF_X1 U627 ( .A(n526), .Z(n527) );
  INV_X1 U628 ( .A(n527), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n528), .A2(n561), .ZN(n578) );
  XNOR2_X1 U630 ( .A(n578), .B(G140), .ZN(G42) );
  XNOR2_X1 U631 ( .A(G116), .B(KEYINPUT117), .ZN(n536) );
  INV_X1 U632 ( .A(n704), .ZN(n531) );
  NOR2_X1 U633 ( .A1(n531), .A2(n366), .ZN(n532) );
  XNOR2_X1 U634 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n533) );
  NAND2_X1 U635 ( .A1(n534), .A2(n543), .ZN(n749) );
  INV_X1 U636 ( .A(n749), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n759), .A2(n576), .ZN(n535) );
  XOR2_X1 U638 ( .A(n536), .B(n535), .Z(G18) );
  INV_X1 U639 ( .A(n724), .ZN(n567) );
  NOR2_X1 U640 ( .A1(n567), .A2(n711), .ZN(n540) );
  XNOR2_X1 U641 ( .A(n540), .B(KEYINPUT30), .ZN(n541) );
  NAND2_X1 U642 ( .A1(n542), .A2(n541), .ZN(n562) );
  NOR2_X1 U643 ( .A1(n544), .A2(n543), .ZN(n599) );
  NAND2_X1 U644 ( .A1(n599), .A2(n527), .ZN(n545) );
  OR2_X1 U645 ( .A1(n562), .A2(n545), .ZN(n756) );
  XNOR2_X1 U646 ( .A(n546), .B(KEYINPUT85), .ZN(n556) );
  INV_X1 U647 ( .A(n711), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n547), .A2(n707), .ZN(n548) );
  NOR2_X1 U649 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U650 ( .A(KEYINPUT28), .B(n550), .Z(n552) );
  NOR2_X1 U651 ( .A1(n552), .A2(n551), .ZN(n570) );
  BUF_X1 U652 ( .A(n553), .Z(n554) );
  NAND2_X1 U653 ( .A1(n570), .A2(n554), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n557), .A2(KEYINPUT47), .ZN(n555) );
  NOR2_X1 U655 ( .A1(n557), .A2(n747), .ZN(n757) );
  NOR2_X1 U656 ( .A1(n557), .A2(n749), .ZN(n754) );
  NOR2_X1 U657 ( .A1(n757), .A2(n754), .ZN(n558) );
  NOR2_X1 U658 ( .A1(KEYINPUT47), .A2(n558), .ZN(n559) );
  XNOR2_X1 U659 ( .A(KEYINPUT38), .B(KEYINPUT79), .ZN(n560) );
  NOR2_X1 U660 ( .A1(n562), .A2(n726), .ZN(n564) );
  XNOR2_X1 U661 ( .A(KEYINPUT77), .B(KEYINPUT39), .ZN(n563) );
  XNOR2_X1 U662 ( .A(n564), .B(n563), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n577), .A2(n758), .ZN(n566) );
  INV_X1 U664 ( .A(n726), .ZN(n720) );
  NOR2_X1 U665 ( .A1(n721), .A2(n567), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n720), .A2(n568), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n569), .B(KEYINPUT41), .ZN(n738) );
  NAND2_X1 U668 ( .A1(n570), .A2(n738), .ZN(n571) );
  BUF_X1 U669 ( .A(n573), .Z(n574) );
  NAND2_X1 U670 ( .A1(n577), .A2(n576), .ZN(n765) );
  XNOR2_X1 U671 ( .A(n580), .B(n579), .ZN(n582) );
  XNOR2_X1 U672 ( .A(n636), .B(n582), .ZN(n581) );
  NAND2_X1 U673 ( .A1(n581), .A2(n369), .ZN(n587) );
  XOR2_X1 U674 ( .A(G227), .B(n582), .Z(n583) );
  NAND2_X1 U675 ( .A1(n583), .A2(G900), .ZN(n584) );
  XNOR2_X1 U676 ( .A(n584), .B(KEYINPUT126), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n585), .A2(G953), .ZN(n586) );
  NAND2_X1 U678 ( .A1(n587), .A2(n586), .ZN(G72) );
  XNOR2_X1 U679 ( .A(n401), .B(G119), .ZN(G21) );
  NAND2_X1 U680 ( .A1(n590), .A2(n366), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n591), .A2(n708), .ZN(n593) );
  XNOR2_X2 U682 ( .A(n595), .B(KEYINPUT91), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT90), .ZN(n603) );
  XNOR2_X1 U684 ( .A(KEYINPUT111), .B(KEYINPUT33), .ZN(n597) );
  XNOR2_X1 U685 ( .A(n598), .B(KEYINPUT34), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n602) );
  XOR2_X1 U687 ( .A(KEYINPUT88), .B(KEYINPUT35), .Z(n601) );
  NOR2_X1 U688 ( .A1(n606), .A2(KEYINPUT44), .ZN(n605) );
  INV_X1 U689 ( .A(KEYINPUT76), .ZN(n604) );
  NOR2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n606), .A2(KEYINPUT76), .ZN(n607) );
  INV_X1 U692 ( .A(n609), .ZN(n621) );
  AND2_X1 U693 ( .A1(n621), .A2(KEYINPUT44), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n610), .A2(KEYINPUT66), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n611), .A2(n366), .ZN(n612) );
  NOR2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n746) );
  XNOR2_X1 U697 ( .A(n614), .B(KEYINPUT104), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT109), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n621), .A2(KEYINPUT66), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n686), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n624), .A2(KEYINPUT44), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  BUF_X1 U705 ( .A(n634), .Z(n635) );
  INV_X1 U706 ( .A(n636), .ZN(n637) );
  BUF_X1 U707 ( .A(n678), .Z(n638) );
  INV_X1 U708 ( .A(n638), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n639), .A2(G478), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(n645) );
  INV_X1 U711 ( .A(n369), .ZN(n644) );
  INV_X1 U712 ( .A(G952), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n683) );
  INV_X1 U714 ( .A(n683), .ZN(n649) );
  NOR2_X1 U715 ( .A1(n645), .A2(n649), .ZN(G63) );
  OR2_X1 U716 ( .A1(n678), .A2(n646), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n650), .A2(n649), .ZN(G66) );
  NOR2_X1 U719 ( .A1(n678), .A2(n651), .ZN(n655) );
  XOR2_X1 U720 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n656), .A2(n683), .ZN(n658) );
  XOR2_X1 U724 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n657) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(G57) );
  INV_X1 U726 ( .A(G210), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n678), .A2(n659), .ZN(n665) );
  XOR2_X1 U728 ( .A(KEYINPUT92), .B(KEYINPUT54), .Z(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT55), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n666), .A2(n683), .ZN(n668) );
  XNOR2_X1 U733 ( .A(KEYINPUT89), .B(KEYINPUT56), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n668), .B(n667), .ZN(G51) );
  INV_X1 U735 ( .A(G475), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n678), .A2(n669), .ZN(n673) );
  XNOR2_X1 U737 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n674), .A2(n683), .ZN(n676) );
  INV_X1 U741 ( .A(KEYINPUT60), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n676), .B(n675), .ZN(G60) );
  INV_X1 U743 ( .A(G469), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n682), .B(n681), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U750 ( .A(n686), .B(G122), .ZN(G24) );
  NOR2_X1 U751 ( .A1(n393), .A2(G953), .ZN(n691) );
  NAND2_X1 U752 ( .A1(G953), .A2(G224), .ZN(n687) );
  XNOR2_X1 U753 ( .A(KEYINPUT61), .B(n687), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n688), .A2(G898), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT123), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n699) );
  XOR2_X1 U757 ( .A(n692), .B(n693), .Z(n695) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U759 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n699), .B(n698), .ZN(G69) );
  NOR2_X1 U762 ( .A1(n700), .A2(KEYINPUT2), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT84), .B(n701), .Z(n703) );
  NAND2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n743) );
  NOR2_X1 U765 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n706), .B(KEYINPUT50), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U768 ( .A(KEYINPUT49), .B(n709), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n366), .A2(n710), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U772 ( .A(KEYINPUT51), .B(n716), .Z(n717) );
  XOR2_X1 U773 ( .A(KEYINPUT119), .B(n717), .Z(n719) );
  INV_X1 U774 ( .A(n738), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n732) );
  NOR2_X1 U776 ( .A1(n720), .A2(n724), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n729) );
  INV_X1 U778 ( .A(n723), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n725), .A2(n724), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U782 ( .A1(n730), .A2(n736), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT52), .ZN(n735) );
  NOR2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n741) );
  INV_X1 U786 ( .A(n736), .ZN(n737) );
  NAND2_X1 U787 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(n449), .ZN(n740) );
  NOR2_X1 U789 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n745) );
  XOR2_X1 U791 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n744) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(G75) );
  INV_X1 U793 ( .A(n746), .ZN(n750) );
  NOR2_X1 U794 ( .A1(n750), .A2(n747), .ZN(n748) );
  XOR2_X1 U795 ( .A(G104), .B(n748), .Z(G6) );
  NOR2_X1 U796 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U799 ( .A(G107), .B(n753), .ZN(G9) );
  XNOR2_X1 U800 ( .A(G128), .B(n754), .ZN(n755) );
  XNOR2_X1 U801 ( .A(n755), .B(KEYINPUT29), .ZN(G30) );
  XNOR2_X1 U802 ( .A(G143), .B(n756), .ZN(G45) );
  XOR2_X1 U803 ( .A(n368), .B(n757), .Z(G48) );
  NAND2_X1 U804 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U805 ( .A(n760), .B(KEYINPUT116), .ZN(n761) );
  XNOR2_X1 U806 ( .A(G113), .B(n761), .ZN(G15) );
  XNOR2_X1 U807 ( .A(n762), .B(KEYINPUT37), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n763), .B(KEYINPUT118), .ZN(n764) );
  XNOR2_X1 U809 ( .A(G125), .B(n764), .ZN(G27) );
  XNOR2_X1 U810 ( .A(G134), .B(n765), .ZN(G36) );
  XOR2_X1 U811 ( .A(G131), .B(n766), .Z(G33) );
  XOR2_X1 U812 ( .A(G137), .B(n767), .Z(G39) );
endmodule

