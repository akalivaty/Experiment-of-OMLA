

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n337), .B(n336), .ZN(n341) );
  XNOR2_X1 U323 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U324 ( .A(n383), .B(KEYINPUT110), .ZN(n384) );
  XNOR2_X1 U325 ( .A(n385), .B(n384), .ZN(n391) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n393), .B(n392), .ZN(n521) );
  XNOR2_X1 U328 ( .A(n342), .B(KEYINPUT64), .ZN(n343) );
  XNOR2_X1 U329 ( .A(n573), .B(n343), .ZN(n555) );
  XNOR2_X1 U330 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n291) );
  XNOR2_X1 U333 ( .A(G99GAT), .B(KEYINPUT83), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U335 ( .A(n292), .B(G190GAT), .Z(n294) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G127GAT), .Z(n368) );
  XNOR2_X1 U337 ( .A(G43GAT), .B(n368), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n299) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n331) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n295), .B(KEYINPUT0), .ZN(n416) );
  XOR2_X1 U342 ( .A(n331), .B(n416), .Z(n297) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U346 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n301) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U349 ( .A(G169GAT), .B(n302), .Z(n404) );
  XOR2_X1 U350 ( .A(G176GAT), .B(G183GAT), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT81), .B(KEYINPUT65), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n404), .B(n305), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n522) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G36GAT), .Z(n309) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G22GAT), .Z(n440) );
  XOR2_X1 U357 ( .A(G1GAT), .B(KEYINPUT71), .Z(n374) );
  XNOR2_X1 U358 ( .A(n440), .B(n374), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U360 ( .A(n310), .B(G197GAT), .Z(n317) );
  XOR2_X1 U361 ( .A(G29GAT), .B(G43GAT), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n358) );
  XOR2_X1 U364 ( .A(n358), .B(KEYINPUT70), .Z(n314) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(n315), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT29), .B(G8GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G15GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U372 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n321) );
  XNOR2_X1 U373 ( .A(KEYINPUT68), .B(KEYINPUT72), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n323), .B(n322), .Z(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n570) );
  XNOR2_X1 U377 ( .A(G176GAT), .B(G92GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(G64GAT), .ZN(n401) );
  XOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .Z(n345) );
  XOR2_X1 U380 ( .A(n401), .B(n345), .Z(n328) );
  NAND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n330) );
  INV_X1 U383 ( .A(KEYINPUT33), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n331), .B(G204GAT), .ZN(n335) );
  XOR2_X1 U386 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n333) );
  XNOR2_X1 U387 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n338), .B(G148GAT), .ZN(n432) );
  XNOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n339), .B(KEYINPUT13), .ZN(n363) );
  XOR2_X1 U393 ( .A(n432), .B(n363), .Z(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n573) );
  INV_X1 U395 ( .A(KEYINPUT41), .ZN(n342) );
  NAND2_X1 U396 ( .A1(n570), .A2(n555), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n344), .B(KEYINPUT46), .ZN(n382) );
  XOR2_X1 U398 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XOR2_X1 U399 ( .A(n398), .B(n345), .Z(n347) );
  NAND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT67), .Z(n349) );
  XNOR2_X1 U403 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U406 ( .A(G50GAT), .B(G162GAT), .Z(n439) );
  XOR2_X1 U407 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n353) );
  XNOR2_X1 U408 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n439), .B(n354), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n357), .B(G92GAT), .Z(n360) );
  XNOR2_X1 U413 ( .A(n358), .B(G106GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n549) );
  XOR2_X1 U415 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n366) );
  XOR2_X1 U416 ( .A(G64GAT), .B(KEYINPUT12), .Z(n362) );
  XNOR2_X1 U417 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n380) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT77), .ZN(n403) );
  XOR2_X1 U423 ( .A(n368), .B(n403), .Z(n370) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT79), .B(G78GAT), .Z(n372) );
  XNOR2_X1 U427 ( .A(G71GAT), .B(G211GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n373), .B(G155GAT), .Z(n376) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U432 ( .A(n378), .B(n377), .Z(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n547) );
  INV_X1 U434 ( .A(n547), .ZN(n577) );
  NOR2_X1 U435 ( .A1(n549), .A2(n577), .ZN(n381) );
  AND2_X1 U436 ( .A1(n382), .A2(n381), .ZN(n385) );
  INV_X1 U437 ( .A(KEYINPUT47), .ZN(n383) );
  XNOR2_X1 U438 ( .A(KEYINPUT36), .B(n549), .ZN(n580) );
  NAND2_X1 U439 ( .A1(n580), .A2(n577), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT111), .ZN(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(n387), .ZN(n388) );
  INV_X1 U442 ( .A(n570), .ZN(n540) );
  NAND2_X1 U443 ( .A1(n388), .A2(n540), .ZN(n389) );
  NOR2_X1 U444 ( .A1(n389), .A2(n573), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n391), .A2(n390), .ZN(n393) );
  XNOR2_X1 U446 ( .A(G211GAT), .B(G218GAT), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n394), .B(KEYINPUT88), .ZN(n395) );
  XOR2_X1 U448 ( .A(n395), .B(KEYINPUT21), .Z(n397) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G204GAT), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n444) );
  XOR2_X1 U451 ( .A(n398), .B(n444), .Z(n400) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U454 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n406), .B(n405), .ZN(n513) );
  NOR2_X1 U457 ( .A1(n521), .A2(n513), .ZN(n407) );
  XNOR2_X1 U458 ( .A(n407), .B(KEYINPUT54), .ZN(n567) );
  XOR2_X1 U459 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n409) );
  XNOR2_X1 U460 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n427) );
  XOR2_X1 U462 ( .A(G162GAT), .B(G148GAT), .Z(n411) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n413) );
  XNOR2_X1 U466 ( .A(G127GAT), .B(G57GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U469 ( .A(G85GAT), .B(n416), .Z(n418) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U474 ( .A(n422), .B(KEYINPUT90), .Z(n425) );
  XNOR2_X1 U475 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(n431), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n566) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n429) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U483 ( .A(n430), .B(KEYINPUT22), .Z(n434) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U486 ( .A(KEYINPUT89), .B(KEYINPUT85), .Z(n436) );
  XNOR2_X1 U487 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U489 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U492 ( .A(n444), .B(n443), .ZN(n460) );
  INV_X1 U493 ( .A(n460), .ZN(n445) );
  AND2_X1 U494 ( .A1(n566), .A2(n445), .ZN(n446) );
  AND2_X1 U495 ( .A1(n567), .A2(n446), .ZN(n447) );
  XNOR2_X1 U496 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U497 ( .A1(n522), .A2(n448), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT119), .B(n449), .Z(n562) );
  NAND2_X1 U499 ( .A1(n562), .A2(n549), .ZN(n452) );
  XOR2_X1 U500 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n450) );
  NOR2_X1 U501 ( .A1(n540), .A2(n573), .ZN(n486) );
  NOR2_X1 U502 ( .A1(n549), .A2(n547), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U504 ( .A(KEYINPUT28), .B(n460), .ZN(n526) );
  XNOR2_X1 U505 ( .A(n513), .B(KEYINPUT27), .ZN(n462) );
  NOR2_X1 U506 ( .A1(n462), .A2(n566), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT93), .ZN(n520) );
  NOR2_X1 U508 ( .A1(n526), .A2(n520), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n522), .A2(n455), .ZN(n469) );
  NOR2_X1 U510 ( .A1(n522), .A2(n513), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n460), .A2(n456), .ZN(n459) );
  XNOR2_X1 U512 ( .A(KEYINPUT25), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT95), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n460), .A2(n522), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U517 ( .A1(n569), .A2(n462), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT94), .B(n463), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT97), .B(n466), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n467), .A2(n566), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n469), .A2(n468), .ZN(n483) );
  NAND2_X1 U523 ( .A1(n470), .A2(n483), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT98), .B(n471), .Z(n498) );
  NAND2_X1 U525 ( .A1(n486), .A2(n498), .ZN(n480) );
  NOR2_X1 U526 ( .A1(n566), .A2(n480), .ZN(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n513), .A2(n480), .ZN(n476) );
  XNOR2_X1 U531 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  NOR2_X1 U534 ( .A1(n522), .A2(n480), .ZN(n479) );
  XNOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  INV_X1 U537 ( .A(n526), .ZN(n517) );
  NOR2_X1 U538 ( .A1(n517), .A2(n480), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NAND2_X1 U541 ( .A1(n580), .A2(n483), .ZN(n484) );
  NOR2_X1 U542 ( .A1(n577), .A2(n484), .ZN(n485) );
  XOR2_X1 U543 ( .A(KEYINPUT37), .B(n485), .Z(n510) );
  NAND2_X1 U544 ( .A1(n486), .A2(n510), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT38), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n496), .A2(n566), .ZN(n489) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n513), .A2(n496), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n522), .A2(n496), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n517), .ZN(n497) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  INV_X1 U559 ( .A(n555), .ZN(n543) );
  NOR2_X1 U560 ( .A1(n543), .A2(n570), .ZN(n509) );
  NAND2_X1 U561 ( .A1(n509), .A2(n498), .ZN(n505) );
  NOR2_X1 U562 ( .A1(n566), .A2(n505), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n501), .Z(G1332GAT) );
  NOR2_X1 U566 ( .A1(n513), .A2(n505), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n522), .A2(n505), .ZN(n504) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n566), .A2(n516), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n516), .ZN(n514) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n522), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  XOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT115), .Z(n529) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n539) );
  INV_X1 U588 ( .A(n522), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n539), .A2(n523), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(n524), .Z(n525) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(KEYINPUT114), .B(n527), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n534), .A2(n570), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n534), .A2(n555), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n577), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n549), .A2(n534), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n537), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n569), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n540), .A2(n550), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n550), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n550), .ZN(n548) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  INV_X1 U616 ( .A(n549), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n552), .Z(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT118), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n570), .A2(n562), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n562), .A2(n555), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT120), .Z(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n577), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT124), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(n565), .Z(n572) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

