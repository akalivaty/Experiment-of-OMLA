//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT3), .A2(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT3), .A2(G107), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(G104), .B2(new_n191), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT3), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(G104), .B2(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n209), .B2(G119), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G119), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(new_n210), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT5), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n212), .A3(G116), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n218));
  OAI211_X1 g032(.A(G113), .B(new_n217), .C1(new_n218), .C2(new_n216), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n206), .A2(KEYINPUT80), .A3(new_n215), .A4(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n215), .A3(new_n200), .A4(new_n204), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n192), .A2(new_n198), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  AND4_X1   g041(.A1(KEYINPUT77), .A2(new_n226), .A3(new_n227), .A4(G101), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n199), .B1(new_n192), .B2(new_n198), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT77), .B1(new_n229), .B2(new_n227), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n207), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n229), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n225), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n237));
  INV_X1    g051(.A(new_n229), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n237), .A2(new_n238), .B1(new_n232), .B2(new_n215), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n227), .A3(G101), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT77), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(KEYINPUT77), .A3(new_n227), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n244), .A3(KEYINPUT79), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n224), .B1(new_n236), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n189), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n224), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n231), .A2(new_n235), .A3(new_n225), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT79), .B1(new_n239), .B2(new_n244), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  OAI211_X1 g074(.A(G128), .B(new_n257), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n262), .B(new_n263), .C1(KEYINPUT1), .C2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT0), .A3(G128), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  MUX2_X1   g085(.A(new_n266), .B(new_n271), .S(G125), .Z(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G224), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n252), .A2(new_n189), .A3(new_n253), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n255), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT81), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n255), .A2(new_n279), .A3(new_n275), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT82), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n221), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n219), .A2(new_n215), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n205), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n283), .A3(new_n205), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n247), .B(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT83), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n272), .B(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(new_n252), .B2(new_n253), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n282), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n281), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n281), .A2(new_n299), .A3(new_n297), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n188), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n264), .A2(G143), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n307), .A2(KEYINPUT96), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(KEYINPUT96), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n264), .A2(G143), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G134), .ZN(new_n313));
  INV_X1    g127(.A(new_n306), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n314), .A2(new_n311), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(KEYINPUT95), .A2(G122), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT95), .A2(G122), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n209), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G122), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G116), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n201), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n201), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n313), .B(new_n317), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n315), .B(new_n316), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n322), .B(KEYINPUT14), .Z(new_n329));
  OAI21_X1  g143(.A(G107), .B1(new_n329), .B2(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT9), .B(G234), .ZN(new_n333));
  INV_X1    g147(.A(G217), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n333), .A2(new_n334), .A3(G953), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n327), .A2(new_n331), .A3(new_n335), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n305), .B1(new_n339), .B2(G902), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  INV_X1    g155(.A(new_n305), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n282), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n343), .A3(KEYINPUT97), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n341), .B2(new_n282), .ZN(new_n346));
  AOI211_X1 g160(.A(G902), .B(new_n305), .C1(new_n337), .C2(new_n338), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G952), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(G234), .A2(G237), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT21), .B(G898), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(G902), .A3(G953), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n344), .A2(new_n348), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G237), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n358), .A2(new_n273), .A3(G143), .A4(G214), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT85), .ZN(new_n360));
  NOR2_X1   g174(.A1(G237), .A2(G953), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G143), .A4(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(G214), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT84), .A3(new_n256), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT84), .B1(new_n365), .B2(new_n256), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT89), .A3(G131), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n372));
  INV_X1    g186(.A(G214), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(G237), .A3(G953), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n374), .B2(G143), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n375), .A2(new_n366), .B1(new_n360), .B2(new_n363), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n370), .A2(new_n378), .A3(new_n379), .A4(KEYINPUT17), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n388), .A2(new_n259), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n259), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n392));
  INV_X1    g206(.A(new_n390), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n388), .A2(new_n259), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n380), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n370), .A2(new_n378), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT93), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n364), .B(new_n377), .C1(new_n367), .C2(new_n368), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT89), .B1(new_n369), .B2(G131), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n376), .A2(new_n371), .A3(new_n377), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n398), .B(new_n400), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT94), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n397), .A2(new_n405), .A3(new_n398), .A4(new_n400), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n396), .A2(new_n399), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n400), .B(KEYINPUT87), .C1(new_n369), .C2(KEYINPUT18), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n376), .B(new_n409), .C1(new_n410), .C2(new_n377), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n376), .A2(new_n377), .ZN(new_n413));
  INV_X1    g227(.A(new_n387), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n259), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(KEYINPUT86), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n387), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(G146), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n413), .A2(KEYINPUT18), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n412), .A2(KEYINPUT88), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(new_n194), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n407), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n282), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G475), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n416), .A2(KEYINPUT19), .A3(new_n418), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n387), .B2(KEYINPUT19), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n434), .A2(new_n436), .A3(new_n259), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n389), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT91), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n397), .A2(new_n400), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(new_n389), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n412), .A2(KEYINPUT88), .A3(new_n420), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT88), .B1(new_n412), .B2(new_n420), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n427), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n428), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n433), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n452), .ZN(new_n454));
  AOI211_X1 g268(.A(KEYINPUT20), .B(new_n454), .C1(new_n428), .C2(new_n450), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n357), .B(new_n432), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G221), .B1(new_n333), .B2(G902), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT75), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n266), .A2(new_n200), .A3(new_n204), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n261), .A2(new_n265), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n205), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .A3(G134), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n316), .A2(G137), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(G134), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI211_X1 g285(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n464), .C2(G134), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT65), .A2(G131), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n470), .B1(new_n316), .B2(G137), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT64), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n468), .A3(new_n470), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n463), .A2(KEYINPUT12), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n463), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT78), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G140), .ZN(new_n488));
  INV_X1    g302(.A(G227), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G953), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n488), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n460), .A2(KEYINPUT10), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n206), .A2(new_n493), .A3(new_n266), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n270), .B1(new_n237), .B2(new_n238), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n492), .A2(new_n494), .B1(new_n495), .B2(new_n244), .ZN(new_n496));
  INV_X1    g310(.A(new_n483), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n486), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n484), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n487), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n492), .A2(new_n494), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(new_n244), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n503), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(G469), .B(G902), .C1(new_n502), .C2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n498), .B1(new_n497), .B2(new_n496), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n485), .A2(new_n486), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n491), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n511), .A3(G469), .ZN(new_n512));
  NAND2_X1  g326(.A1(G469), .A2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n459), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n456), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G472), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n270), .B1(new_n476), .B2(new_n482), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n469), .A2(new_n466), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n261), .A2(new_n521), .A3(new_n265), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n377), .B2(new_n481), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n233), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n475), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n479), .A2(new_n480), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n474), .B1(new_n526), .B2(new_n467), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n271), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n233), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n266), .B(new_n521), .C1(G131), .C2(new_n473), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n518), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n361), .A2(G210), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT68), .Z(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n536), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n533), .A2(new_n534), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n282), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n524), .A2(new_n531), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n540), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n534), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n519), .A2(new_n523), .A3(new_n233), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT30), .B1(new_n519), .B2(new_n523), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n528), .A2(new_n552), .A3(new_n530), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n554), .B2(new_n233), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n549), .B(new_n541), .C1(new_n548), .C2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n544), .B1(new_n556), .B2(KEYINPUT72), .ZN(new_n557));
  INV_X1    g371(.A(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n540), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n541), .A4(new_n549), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n517), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n555), .B2(new_n548), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n529), .B1(new_n551), .B2(new_n553), .ZN(new_n566));
  NOR4_X1   g380(.A1(new_n566), .A2(KEYINPUT69), .A3(new_n540), .A4(new_n550), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n546), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n524), .B2(new_n531), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n540), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n555), .A2(new_n568), .A3(new_n548), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT71), .B(new_n540), .C1(new_n571), .C2(new_n572), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n563), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT32), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n563), .C1(new_n569), .C2(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n562), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n334), .B1(G234), .B2(new_n282), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n212), .B2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n264), .A2(KEYINPUT23), .A3(G119), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n587), .B(new_n588), .C1(G119), .C2(new_n264), .ZN(new_n589));
  XNOR2_X1  g403(.A(G119), .B(G128), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT24), .B(G110), .Z(new_n591));
  OAI22_X1  g405(.A1(new_n589), .A2(G110), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n389), .A2(new_n592), .A3(new_n415), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n393), .B2(new_n394), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(G110), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT73), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n593), .B(new_n601), .C1(new_n595), .C2(new_n597), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n282), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n603), .A2(KEYINPUT25), .A3(new_n282), .A4(new_n604), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n585), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n603), .A2(new_n604), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n585), .A2(new_n282), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT74), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n583), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n303), .A2(new_n516), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  OAI21_X1  g432(.A(new_n282), .B1(new_n569), .B2(new_n578), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n579), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n614), .B(new_n459), .C1(new_n508), .C2(new_n514), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  INV_X1    g441(.A(new_n430), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n628), .B2(new_n428), .ZN(new_n629));
  INV_X1    g443(.A(G475), .ZN(new_n630));
  OAI22_X1  g444(.A1(new_n453), .A2(new_n455), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n341), .A2(new_n304), .A3(new_n282), .ZN(new_n632));
  NAND2_X1  g446(.A1(G478), .A2(G902), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n332), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n341), .B(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n632), .B(new_n633), .C1(new_n637), .C2(new_n304), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n631), .A2(new_n356), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n303), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n627), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n344), .A2(new_n348), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n356), .B(KEYINPUT100), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n631), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT101), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(KEYINPUT101), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n303), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n627), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n598), .B(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n612), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n609), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n620), .A2(new_n579), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n620), .A2(new_n663), .A3(new_n579), .A4(new_n660), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n303), .A2(new_n516), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  OR2_X1    g481(.A1(new_n355), .A2(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n352), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n631), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n303), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n583), .A2(new_n515), .A3(new_n659), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n264), .ZN(G30));
  AOI21_X1  g490(.A(new_n299), .B1(new_n281), .B2(new_n297), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n300), .B(new_n296), .C1(new_n278), .C2(new_n280), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT38), .Z(new_n680));
  INV_X1    g494(.A(new_n515), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n669), .B(KEYINPUT39), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n187), .B(new_n659), .C1(new_n683), .C2(KEYINPUT40), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(KEYINPUT40), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n631), .A2(new_n645), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n580), .A2(new_n582), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n567), .B(new_n565), .C1(new_n540), .C2(new_n545), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n680), .A2(new_n685), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT103), .B(G143), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  NAND3_X1  g508(.A1(new_n631), .A2(new_n639), .A3(new_n669), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n303), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n674), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT104), .B(G146), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G48));
  INV_X1    g514(.A(G469), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n502), .A2(new_n507), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n702), .B2(new_n282), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n508), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n459), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n583), .A2(new_n615), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n303), .A3(new_n640), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n650), .A2(new_n303), .A3(new_n651), .A4(new_n706), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT105), .B(G116), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  NOR2_X1   g526(.A1(new_n583), .A2(new_n659), .ZN(new_n713));
  INV_X1    g527(.A(new_n456), .ZN(new_n714));
  INV_X1    g528(.A(new_n705), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n303), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR3_X1   g531(.A1(new_n519), .A2(new_n523), .A3(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n552), .B1(new_n528), .B2(new_n530), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n233), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n548), .A3(new_n531), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT69), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n555), .A2(new_n564), .A3(new_n548), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n533), .A2(new_n725), .A3(new_n534), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n532), .B2(new_n572), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n540), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(KEYINPUT107), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n576), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT107), .B1(new_n724), .B2(new_n728), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n563), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n703), .A2(new_n508), .A3(new_n458), .A4(new_n648), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n614), .A2(new_n732), .A3(new_n620), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n303), .A3(new_n687), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT108), .B(G122), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G24));
  AND3_X1   g551(.A1(new_n732), .A2(new_n620), .A3(new_n660), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n303), .A2(new_n738), .A3(new_n696), .A4(new_n715), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NOR3_X1   g554(.A1(new_n677), .A2(new_n678), .A3(new_n188), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n513), .B(KEYINPUT109), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n512), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n702), .A2(new_n701), .A3(new_n282), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n458), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n631), .A2(new_n639), .A3(new_n669), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n616), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n741), .A2(new_n616), .A3(new_n746), .A4(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  AND2_X1   g566(.A1(new_n741), .A2(new_n616), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n671), .A2(new_n745), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  OR2_X1    g570(.A1(new_n631), .A2(new_n638), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT43), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT110), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n624), .A3(new_n660), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n509), .A2(new_n511), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n701), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT46), .B1(new_n766), .B2(new_n742), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n508), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n458), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n682), .A3(new_n741), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n760), .B2(new_n761), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  XOR2_X1   g588(.A(new_n770), .B(KEYINPUT47), .Z(new_n775));
  INV_X1    g589(.A(new_n741), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n696), .A2(new_n583), .A3(new_n615), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n382), .ZN(G42));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n758), .A2(new_n352), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n732), .A2(new_n620), .A3(new_n614), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n741), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n704), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n775), .B1(new_n459), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n783), .B2(KEYINPUT112), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n776), .A2(new_n705), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(new_n738), .A3(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n691), .A2(new_n615), .A3(new_n352), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n631), .A2(new_n639), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n781), .A2(new_n782), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n705), .A2(new_n187), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT114), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n680), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n796), .A2(KEYINPUT50), .A3(new_n799), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n789), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n785), .A2(new_n788), .A3(KEYINPUT113), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n780), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT115), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n631), .A2(new_n639), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n340), .A2(new_n343), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n631), .B2(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n621), .A2(new_n625), .A3(new_n622), .A4(new_n648), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n303), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n716), .A2(new_n707), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n665), .A2(new_n735), .A3(new_n617), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n710), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n631), .A2(new_n810), .A3(new_n670), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n713), .A2(new_n681), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n738), .A2(new_n746), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n741), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n751), .A2(new_n821), .A3(new_n755), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n715), .B(new_n187), .C1(new_n677), .C2(new_n678), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n695), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n187), .B1(new_n677), .B2(new_n678), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n686), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n745), .A2(new_n659), .A3(new_n669), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n688), .B2(new_n690), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n826), .A2(new_n738), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n673), .B(new_n303), .C1(new_n671), .C2(new_n696), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n824), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n303), .A2(new_n830), .A3(new_n687), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n824), .A2(new_n832), .A3(new_n739), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT111), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n832), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n739), .A2(new_n834), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT52), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n831), .A2(new_n824), .A3(new_n832), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n823), .A2(new_n836), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n833), .A2(new_n835), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n823), .A2(new_n847), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(KEYINPUT53), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n852), .B2(KEYINPUT54), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n785), .B2(new_n788), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(new_n804), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n855), .B2(new_n804), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n781), .A2(new_n616), .A3(new_n790), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(KEYINPUT48), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(KEYINPUT48), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n796), .A2(new_n303), .A3(new_n715), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n350), .C1(new_n809), .C2(new_n793), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n862), .B(new_n864), .C1(new_n860), .C2(new_n858), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n808), .A2(new_n853), .A3(new_n857), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n349), .A2(new_n273), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n786), .A2(KEYINPUT49), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n786), .A2(KEYINPUT49), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n615), .A2(new_n188), .A3(new_n458), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OR4_X1    g686(.A1(new_n680), .A2(new_n691), .A3(new_n757), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n273), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n845), .A2(new_n848), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(G902), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n255), .A2(new_n276), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n275), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n876), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n880), .B2(new_n883), .ZN(G51));
  NOR2_X1   g699(.A1(new_n878), .A2(new_n766), .ZN(new_n886));
  INV_X1    g700(.A(new_n702), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n742), .B(KEYINPUT118), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT57), .Z(new_n889));
  AOI21_X1  g703(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n849), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n889), .C1(new_n849), .C2(new_n890), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n887), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n893), .B1(new_n900), .B2(new_n889), .ZN(new_n901));
  INV_X1    g715(.A(new_n894), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n702), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n875), .B1(new_n897), .B2(new_n904), .ZN(G54));
  AND3_X1   g719(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n876), .B1(new_n906), .B2(new_n451), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n451), .B2(new_n906), .ZN(G60));
  INV_X1    g722(.A(new_n637), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n633), .B(KEYINPUT59), .Z(new_n910));
  AOI211_X1 g724(.A(new_n909), .B(new_n910), .C1(new_n898), .C2(new_n899), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n853), .A2(new_n910), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n875), .B(new_n911), .C1(new_n912), .C2(new_n909), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  AOI21_X1  g729(.A(new_n610), .B1(new_n877), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n875), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n917), .B2(KEYINPUT121), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n877), .A2(new_n657), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G66));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n353), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n817), .B(KEYINPUT122), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n925), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n881), .B1(G898), .B2(new_n273), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT123), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  NAND3_X1  g743(.A1(new_n434), .A2(new_n438), .A3(new_n436), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT124), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n554), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n778), .B1(new_n762), .B2(new_n772), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n832), .A2(new_n739), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT125), .Z(new_n935));
  NAND4_X1  g749(.A1(new_n828), .A2(new_n770), .A3(new_n616), .A4(new_n682), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n751), .A2(new_n755), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT127), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n933), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n273), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n489), .A2(G900), .A3(G953), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n932), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n812), .B(KEYINPUT126), .Z(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n681), .A3(new_n682), .A4(new_n753), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n935), .A2(new_n692), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n933), .B(new_n945), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n273), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n942), .B1(new_n952), .B2(new_n932), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n939), .B2(new_n924), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n558), .A2(new_n548), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n875), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n925), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n949), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n548), .A3(new_n558), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n722), .A2(new_n559), .A3(new_n723), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n852), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n961), .A3(new_n963), .ZN(G57));
endmodule


