//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n219), .B1(new_n202), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G77), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n218), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n215), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n216), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n256), .B1(G150), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(KEYINPUT67), .B1(G20), .B2(new_n203), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n249), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n215), .A3(new_n247), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n264), .A2(new_n266), .B1(G50), .B2(new_n263), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(G274), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n277), .B2(new_n220), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n281), .B1(new_n225), .B2(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n268), .B1(new_n269), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G179), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n268), .A2(KEYINPUT9), .B1(new_n287), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n261), .B2(new_n267), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n286), .A2(new_n296), .A3(G190), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(new_n286), .B2(G190), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n292), .A3(new_n303), .A4(new_n294), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n291), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  OAI211_X1 g0108(.A(G232), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n279), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n285), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n272), .A2(G238), .A3(new_n276), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n275), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n306), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT13), .B(new_n318), .C1(new_n315), .C2(new_n285), .ZN(new_n321));
  OAI21_X1  g0121(.A(G169), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n306), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(new_n319), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT72), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n316), .A2(new_n328), .A3(new_n306), .A4(new_n319), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n325), .A2(new_n327), .A3(G179), .A4(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n324), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(KEYINPUT75), .A3(G169), .A4(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(G169), .B(new_n333), .C1(new_n320), .C2(new_n321), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n256), .A2(G77), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n249), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT11), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n263), .A2(G68), .B1(KEYINPUT73), .B2(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n264), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G68), .A3(new_n265), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT15), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G87), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n256), .ZN(new_n359));
  INV_X1    g0159(.A(new_n257), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n251), .A2(new_n253), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n359), .B1(new_n216), .B2(new_n225), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n263), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(new_n248), .B1(new_n225), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n249), .A2(G77), .A3(new_n263), .A4(new_n265), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT68), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n275), .B1(new_n277), .B2(new_n224), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n279), .A2(G232), .A3(new_n280), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n279), .A2(G238), .A3(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n279), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(new_n285), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(KEYINPUT69), .B1(G190), .B2(new_n374), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n352), .B1(new_n332), .B2(G200), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n325), .A2(new_n327), .A3(G190), .A4(new_n329), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n374), .A2(G169), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n289), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n368), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n380), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n254), .A2(new_n265), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n348), .B1(new_n363), .B2(new_n361), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n250), .A2(new_n341), .ZN(new_n391));
  OAI21_X1  g0191(.A(G20), .B1(new_n391), .B2(new_n201), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n257), .A2(G159), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n279), .B2(G20), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n307), .A2(new_n308), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n394), .B1(new_n399), .B2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n249), .B1(new_n400), .B2(KEYINPUT16), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n341), .B1(new_n396), .B2(new_n398), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n390), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n220), .A2(G1698), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G223), .B2(G1698), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n407), .A2(new_n397), .B1(new_n270), .B2(new_n354), .ZN(new_n408));
  INV_X1    g0208(.A(G274), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n285), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n408), .A2(new_n285), .B1(new_n274), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  INV_X1    g0212(.A(G232), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n277), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n272), .A2(KEYINPUT76), .A3(G232), .A4(new_n276), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n269), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n411), .A2(new_n416), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(G179), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT18), .B1(new_n405), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT7), .B1(new_n397), .B2(new_n216), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n307), .A2(new_n308), .A3(new_n395), .A4(G20), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n394), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n404), .A2(new_n426), .A3(new_n248), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(G200), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n411), .A2(new_n416), .A3(G190), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n389), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n375), .B1(new_n411), .B2(new_n416), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n419), .B2(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n405), .A2(new_n434), .A3(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n418), .A2(G169), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n289), .B2(new_n418), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n427), .A2(new_n389), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n421), .A2(new_n432), .A3(new_n435), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n305), .A2(new_n353), .A3(new_n387), .A4(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n216), .B(G87), .C1(new_n307), .C2(new_n308), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT22), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT22), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n279), .A2(new_n446), .A3(new_n216), .A4(G87), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OR3_X1    g0251(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n452));
  OAI211_X1 g0252(.A(KEYINPUT80), .B(KEYINPUT23), .C1(new_n216), .C2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n216), .A2(G33), .A3(G116), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n448), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n451), .A2(new_n453), .A3(new_n452), .A4(new_n454), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n445), .B2(new_n447), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n461), .A3(new_n248), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n263), .A2(G107), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT25), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT77), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n270), .B2(G1), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n262), .A2(KEYINPUT77), .A3(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n264), .A2(new_n469), .A3(new_n372), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT81), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n463), .B(KEYINPUT25), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n264), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G257), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n478));
  OAI211_X1 g0278(.A(G250), .B(new_n280), .C1(new_n307), .C2(new_n308), .ZN(new_n479));
  INV_X1    g0279(.A(G294), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n478), .B(new_n479), .C1(new_n270), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n262), .A2(G45), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n285), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n481), .A2(new_n285), .B1(new_n485), .B2(G264), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n484), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n410), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(G190), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n481), .A2(new_n285), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(G264), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n462), .A2(new_n477), .A3(new_n489), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n484), .A2(new_n483), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G257), .A3(new_n272), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(new_n280), .C1(new_n307), .C2(new_n308), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n285), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n269), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n498), .A2(new_n506), .A3(new_n289), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n205), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n372), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n257), .A2(G77), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n372), .B1(new_n396), .B2(new_n398), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n248), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n263), .A2(G97), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n473), .B2(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n508), .A2(new_n509), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n422), .B2(new_n423), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n249), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n521), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n498), .A2(new_n506), .A3(G190), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n497), .B1(new_n285), .B2(new_n505), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n529), .C1(new_n375), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n494), .A2(new_n523), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n533));
  OAI211_X1 g0333(.A(G238), .B(new_n280), .C1(new_n307), .C2(new_n308), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n534), .C1(new_n270), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n285), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n272), .A2(G274), .A3(new_n483), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n272), .A2(G250), .A3(new_n482), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(G179), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n285), .B2(new_n536), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n269), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n216), .B1(new_n313), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G87), .B2(new_n206), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n216), .B(G68), .C1(new_n307), .C2(new_n308), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n255), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n358), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n551), .A2(new_n248), .B1(new_n363), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n473), .A2(new_n358), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n248), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n363), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n544), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n473), .A2(G87), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n543), .A2(G190), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n537), .A2(new_n541), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n532), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n279), .A2(G264), .A3(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n279), .A2(G257), .A3(new_n280), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n397), .A2(G303), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n285), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n485), .A2(G270), .B1(new_n487), .B2(new_n410), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n473), .A2(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n363), .A2(new_n535), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n535), .A2(G20), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n248), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n503), .B(new_n216), .C1(G33), .C2(new_n549), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND4_X1   g0382(.A1(KEYINPUT20), .A2(new_n581), .A3(new_n248), .A4(new_n579), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n578), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(new_n584), .A3(KEYINPUT21), .A4(G169), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n269), .B1(new_n574), .B2(new_n575), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(KEYINPUT79), .A3(KEYINPUT21), .A4(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n584), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n574), .A2(new_n575), .A3(G179), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n584), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n584), .B1(new_n576), .B2(G200), .ZN(new_n596));
  INV_X1    g0396(.A(G190), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n576), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n590), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n249), .B1(new_n456), .B2(new_n457), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n461), .B1(new_n476), .B2(new_n471), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n492), .A2(new_n269), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n486), .A2(new_n289), .A3(new_n488), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT82), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n492), .A2(G179), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n486), .B2(new_n488), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n248), .B1(new_n460), .B2(KEYINPUT24), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n456), .A2(new_n457), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n477), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT82), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n569), .A2(new_n599), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n443), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT83), .ZN(G372));
  INV_X1    g0417(.A(new_n291), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n421), .A2(new_n440), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n323), .A2(new_n330), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n337), .B2(new_n334), .ZN(new_n621));
  INV_X1    g0421(.A(new_n383), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n621), .A2(new_n351), .B1(new_n622), .B2(new_n386), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n435), .A2(new_n432), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n301), .A2(new_n304), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n618), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n565), .A2(G169), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n542), .B1(new_n553), .B2(new_n555), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n523), .A2(new_n531), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n553), .B(new_n562), .C1(new_n543), .C2(new_n375), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT84), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(G190), .B2(new_n543), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n563), .A2(KEYINPUT84), .A3(new_n566), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(new_n639), .A3(new_n494), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n609), .A2(new_n612), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n590), .A2(new_n641), .A3(new_n595), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n633), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n523), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT26), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n568), .A2(new_n647), .A3(new_n523), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n630), .B1(new_n443), .B2(new_n650), .ZN(G369));
  NAND3_X1  g0451(.A1(new_n262), .A2(new_n216), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n584), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n599), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n590), .A2(new_n595), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT85), .B(G330), .Z(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n605), .B1(new_n601), .B2(new_n604), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n609), .A2(new_n612), .A3(KEYINPUT82), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n666), .A2(new_n667), .A3(new_n494), .ZN(new_n668));
  INV_X1    g0468(.A(new_n657), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n601), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n609), .A2(new_n612), .A3(new_n657), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n641), .A2(new_n657), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n660), .A2(new_n657), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  NOR3_X1   g0477(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n209), .A2(new_n271), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(G1), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n213), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n669), .B1(new_n644), .B2(new_n649), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n647), .B1(new_n568), .B2(new_n523), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n645), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT88), .B(new_n647), .C1(new_n568), .C2(new_n523), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n666), .A2(new_n667), .A3(new_n590), .A4(new_n595), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n633), .B1(new_n693), .B2(new_n640), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT29), .B(new_n669), .C1(new_n691), .C2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n565), .A2(KEYINPUT86), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(new_n507), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n576), .A2(new_n492), .A3(new_n289), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n543), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n698), .A2(new_n700), .A3(KEYINPUT87), .A4(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT87), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n697), .A2(new_n507), .A3(new_n702), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n498), .A2(new_n506), .A3(new_n543), .A4(new_n486), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n593), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n543), .A2(new_n486), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n594), .A2(new_n711), .A3(KEYINPUT30), .A4(new_n530), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n707), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n615), .A2(KEYINPUT31), .B1(new_n657), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n669), .A2(new_n715), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n663), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n696), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n682), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n661), .A2(new_n663), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n216), .A2(G13), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n262), .B1(new_n726), .B2(G45), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n725), .B(new_n665), .C1(new_n679), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n727), .ZN(new_n729));
  INV_X1    g0529(.A(new_n679), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n279), .A2(new_n209), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(G116), .B2(new_n209), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n242), .A2(new_n273), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n397), .A2(new_n209), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n273), .B2(new_n214), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT89), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n215), .B1(G20), .B2(new_n269), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n731), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n597), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n289), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n549), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n216), .A2(new_n289), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n597), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n216), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n202), .B1(new_n758), .B2(new_n354), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(G190), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n752), .B(new_n759), .C1(G68), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n597), .A3(G200), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n279), .B1(new_n762), .B2(new_n372), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT32), .A3(G159), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT32), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n763), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n748), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n761), .B(new_n771), .C1(new_n250), .C2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n764), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT91), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT91), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n225), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n279), .B1(new_n766), .B2(G329), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n758), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n786), .A2(new_n760), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n774), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n784), .B(new_n788), .C1(G322), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n762), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n755), .A2(G326), .B1(new_n791), .B2(G283), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n790), .B(new_n792), .C1(new_n480), .C2(new_n751), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n775), .A2(new_n781), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n747), .B1(new_n796), .B2(new_n744), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n742), .B(KEYINPUT93), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n661), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT94), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n728), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  INV_X1    g0603(.A(new_n731), .ZN(new_n804));
  INV_X1    g0604(.A(new_n649), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n637), .A2(new_n638), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n633), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n532), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n632), .B1(new_n808), .B2(new_n642), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n657), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n386), .A2(new_n657), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n368), .A2(new_n657), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n380), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n813), .B2(new_n386), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n683), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n804), .B1(new_n818), .B2(new_n722), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT96), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n722), .B2(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n762), .A2(new_n354), .ZN(new_n825));
  INV_X1    g0625(.A(new_n760), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n826), .A2(new_n827), .B1(new_n372), .B2(new_n758), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n825), .B(new_n828), .C1(G303), .C2(new_n755), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n397), .B1(new_n765), .B2(new_n794), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n830), .B(new_n752), .C1(G294), .C2(new_n789), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n535), .C2(new_n780), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G137), .A2(new_n755), .B1(new_n760), .B2(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n774), .C1(new_n780), .C2(new_n769), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT95), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT34), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n279), .B1(new_n765), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G68), .B2(new_n791), .ZN(new_n840));
  INV_X1    g0640(.A(new_n758), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G50), .A2(new_n841), .B1(new_n750), .B2(G58), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n836), .A2(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n744), .ZN(new_n846));
  INV_X1    g0646(.A(G77), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n744), .A2(new_n739), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n804), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n846), .B(new_n849), .C1(new_n740), .C2(new_n814), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n824), .A2(new_n850), .ZN(G384));
  OR2_X1    g0651(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n217), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OR3_X1    g0655(.A1(new_n225), .A2(new_n213), .A3(new_n391), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n202), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n262), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n443), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n685), .A2(new_n695), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n685), .A2(new_n695), .A3(new_n860), .A4(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n630), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT104), .Z(new_n867));
  INV_X1    g0667(.A(KEYINPUT97), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n339), .B2(new_n352), .ZN(new_n869));
  AOI211_X1 g0669(.A(KEYINPUT97), .B(new_n351), .C1(new_n331), .C2(new_n338), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n351), .A2(new_n669), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n383), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n621), .B2(new_n383), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT98), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT97), .B1(new_n621), .B2(new_n351), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n339), .A2(new_n868), .A3(new_n352), .ZN(new_n878));
  INV_X1    g0678(.A(new_n873), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT98), .ZN(new_n881));
  INV_X1    g0681(.A(new_n875), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT99), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n403), .B2(new_n394), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n424), .A2(KEYINPUT99), .A3(new_n425), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n402), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n390), .B1(new_n888), .B2(new_n401), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n430), .B1(new_n889), .B2(new_n420), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n655), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n437), .A2(new_n438), .ZN(new_n893));
  INV_X1    g0693(.A(new_n655), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n438), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n430), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n441), .A2(new_n891), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT100), .A4(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n899), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n811), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n815), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n884), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AND4_X1   g0710(.A1(KEYINPUT39), .A2(new_n902), .A3(new_n903), .A4(new_n906), .ZN(new_n911));
  XNOR2_X1  g0711(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n912));
  INV_X1    g0712(.A(new_n895), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n441), .A2(KEYINPUT102), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n893), .A2(new_n895), .A3(new_n430), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n897), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT102), .B1(new_n441), .B2(new_n913), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT39), .B1(new_n920), .B2(new_n900), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n657), .B1(new_n877), .B2(new_n878), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n619), .A2(new_n655), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n910), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n867), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n713), .B1(new_n706), .B2(new_n703), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT106), .B1(new_n929), .B2(new_n719), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n707), .A2(new_n714), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n718), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n814), .B1(new_n935), .B2(new_n717), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n937), .B(new_n907), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n920), .B2(new_n900), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n937), .B(new_n945), .C1(new_n938), .C2(new_n939), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n615), .A2(KEYINPUT31), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n716), .A2(new_n657), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n933), .B2(new_n930), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n443), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n663), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n947), .B2(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n928), .A2(new_n953), .B1(new_n262), .B2(new_n726), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n928), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n859), .B1(new_n954), .B2(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n634), .B1(new_n528), .B2(new_n669), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n523), .B2(new_n669), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT107), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n673), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n613), .B2(new_n606), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n657), .B1(new_n963), .B2(new_n523), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n668), .A3(new_n675), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n563), .A2(new_n669), .ZN(new_n968));
  MUX2_X1   g0768(.A(new_n807), .B(new_n633), .S(new_n968), .Z(new_n969));
  OAI22_X1  g0769(.A1(new_n964), .A2(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n967), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n962), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n961), .B(KEYINPUT108), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n679), .B(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n676), .A2(new_n958), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n676), .A2(new_n958), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n665), .A3(new_n672), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n673), .A3(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n675), .A2(new_n668), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n672), .B2(new_n675), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n665), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n723), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n978), .B1(new_n992), .B2(new_n723), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n977), .B1(new_n993), .B2(new_n729), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n745), .B1(new_n209), .B2(new_n552), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n238), .A2(new_n736), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n731), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G137), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n279), .B1(new_n765), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n751), .A2(new_n341), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G150), .C2(new_n789), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n826), .A2(new_n769), .B1(new_n756), .B2(new_n834), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n250), .A2(new_n758), .B1(new_n762), .B2(new_n225), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(new_n780), .C2(new_n202), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n774), .A2(new_n783), .B1(new_n756), .B2(new_n794), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n780), .A2(new_n827), .B1(KEYINPUT110), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n397), .B1(new_n765), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G97), .B2(new_n791), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n760), .A2(G294), .B1(new_n750), .B2(G107), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n841), .A2(G116), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT46), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1005), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n997), .B1(new_n1017), .B2(new_n744), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n969), .A2(new_n798), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n994), .A2(new_n1020), .ZN(G387));
  OAI22_X1  g0821(.A1(new_n678), .A2(new_n733), .B1(G107), .B2(new_n209), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n235), .A2(new_n273), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  INV_X1    g0824(.A(new_n678), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n1025), .C1(G68), .C2(G77), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n254), .A2(new_n202), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT50), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n736), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1022), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n731), .B1(new_n1030), .B2(new_n746), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n756), .A2(new_n769), .B1(new_n751), .B2(new_n552), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n279), .B1(new_n549), .B2(new_n762), .C1(new_n774), .C2(new_n202), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n254), .C2(new_n760), .ZN(new_n1034));
  INV_X1    g0834(.A(G150), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n758), .A2(new_n225), .B1(new_n765), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT112), .Z(new_n1037));
  OAI211_X1 g0837(.A(new_n1034), .B(new_n1037), .C1(new_n341), .C2(new_n780), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n279), .B1(new_n766), .B2(G326), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n751), .A2(new_n827), .B1(new_n758), .B2(new_n480), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G311), .A2(new_n760), .B1(new_n755), .B2(G322), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n1009), .B2(new_n774), .C1(new_n780), .C2(new_n783), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1039), .B1(new_n535), .B2(new_n762), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1038), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1031), .B1(new_n1049), .B2(new_n744), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n670), .A2(new_n671), .A3(new_n798), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n990), .A2(new_n729), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n991), .A2(new_n730), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n723), .A2(new_n990), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n987), .A2(new_n991), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n992), .A2(new_n730), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n987), .A2(new_n727), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n960), .A2(new_n743), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n745), .B1(new_n549), .B2(new_n209), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n245), .A2(new_n736), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n731), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n841), .A2(G68), .B1(new_n766), .B2(G143), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n826), .A2(new_n202), .B1(new_n751), .B2(new_n847), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n397), .A4(new_n825), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(KEYINPUT113), .B2(new_n1063), .C1(new_n361), .C2(new_n780), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n789), .A2(G159), .B1(G150), .B2(new_n755), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n279), .B1(new_n766), .B2(G322), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n372), .B2(new_n762), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n826), .A2(new_n783), .B1(new_n751), .B2(new_n535), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G283), .C2(new_n841), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n780), .B2(new_n480), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n789), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1067), .A2(new_n1069), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1062), .B1(new_n1077), .B2(new_n744), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1058), .B1(new_n1059), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1057), .A2(new_n1079), .ZN(G390));
  INV_X1    g0880(.A(G330), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n950), .A2(new_n443), .A3(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n629), .B(new_n1082), .C1(new_n863), .C2(new_n864), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n663), .B(new_n814), .C1(new_n717), .C2(new_n721), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n938), .B2(new_n939), .ZN(new_n1086));
  OAI211_X1 g0886(.A(G330), .B(new_n814), .C1(new_n935), .C2(new_n717), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n876), .A2(new_n883), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n632), .B1(new_n808), .B2(new_n692), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n657), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n813), .A2(new_n386), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n811), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1086), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n909), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n950), .A2(new_n1081), .A3(new_n816), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n938), .B2(new_n939), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n876), .A2(new_n883), .A3(new_n1084), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1083), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT114), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1083), .B(new_n1102), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1097), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n909), .B1(new_n938), .B2(new_n939), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n923), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n922), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n920), .A2(new_n900), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1107), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1093), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n884), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1105), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n938), .B2(new_n939), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n923), .B1(new_n884), .B2(new_n909), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1086), .C1(new_n1116), .C2(new_n922), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n730), .B1(new_n1104), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n729), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n756), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n397), .B1(new_n766), .B2(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n826), .B2(new_n998), .C1(new_n838), .C2(new_n774), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n758), .A2(new_n1035), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT53), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n751), .A2(new_n769), .B1(new_n762), .B2(new_n202), .ZN(new_n1130));
  OR4_X1    g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n780), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n780), .A2(new_n549), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n789), .A2(G116), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G68), .A2(new_n791), .B1(new_n750), .B2(G77), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G107), .A2(new_n760), .B1(new_n755), .B2(G283), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n397), .B1(new_n765), .B2(new_n480), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G87), .B2(new_n841), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1131), .A2(new_n1133), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n744), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n804), .B1(new_n361), .B2(new_n848), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n922), .C2(new_n740), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1122), .A2(new_n1123), .A3(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1082), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n865), .A2(new_n630), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT57), .B1(new_n1121), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n936), .B1(new_n876), .B2(new_n883), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n941), .B1(new_n1151), .B2(new_n907), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n946), .A2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n943), .A2(KEYINPUT117), .A3(G330), .A4(new_n946), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n268), .A2(new_n655), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT55), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n305), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1150), .B(new_n1162), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n926), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n927), .A3(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1146), .B1(new_n1149), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1121), .A2(new_n1148), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1169), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n909), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1086), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1102), .B1(new_n1175), .B2(new_n1083), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1103), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1118), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1169), .B1(new_n1178), .B2(new_n1083), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1161), .A2(new_n927), .A3(new_n1163), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n927), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1182), .A3(KEYINPUT118), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1168), .A2(new_n1171), .A3(new_n1183), .A4(new_n730), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1000), .B1(G116), .B2(new_n755), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT115), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n279), .A2(G41), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n827), .B2(new_n765), .C1(new_n225), .C2(new_n758), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n826), .A2(new_n549), .B1(new_n762), .B2(new_n250), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G107), .C2(new_n789), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1186), .B(new_n1190), .C1(new_n552), .C2(new_n780), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1187), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n758), .A2(new_n1132), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n826), .A2(new_n838), .B1(new_n751), .B2(new_n1035), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G125), .C2(new_n755), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n1124), .B2(new_n774), .C1(new_n998), .C2(new_n780), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n791), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1196), .B1(new_n1192), .B2(new_n1191), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n744), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n804), .B1(new_n202), .B2(new_n848), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1162), .C2(new_n740), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1167), .B2(new_n727), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1184), .A2(new_n1211), .ZN(G375));
  NAND3_X1  g1012(.A1(new_n1173), .A2(new_n1148), .A3(new_n1174), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1101), .A2(new_n1103), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(new_n978), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT119), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1175), .A2(new_n729), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n804), .B1(new_n341), .B2(new_n848), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n744), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n279), .B1(new_n765), .B2(new_n1124), .C1(new_n250), .C2(new_n762), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G159), .A2(new_n841), .B1(new_n750), .B2(G50), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n756), .B2(new_n838), .C1(new_n826), .C2(new_n1132), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(G137), .C2(new_n789), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n779), .A2(G150), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n779), .A2(G107), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n279), .B1(new_n766), .B2(G303), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n751), .B2(new_n552), .C1(new_n774), .C2(new_n827), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n826), .A2(new_n535), .B1(new_n549), .B2(new_n758), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n756), .A2(new_n480), .B1(new_n762), .B2(new_n847), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1223), .A2(new_n1224), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1218), .B1(new_n1219), .B2(new_n1231), .C1(new_n884), .C2(new_n740), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1217), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1216), .A2(new_n1234), .ZN(G381));
  AND3_X1   g1035(.A1(new_n1122), .A2(new_n1123), .A3(new_n1144), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n994), .A3(new_n1020), .A4(new_n1237), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1238), .A2(G375), .A3(G381), .ZN(G407));
  NAND2_X1  g1039(.A1(new_n656), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G375), .C2(new_n1242), .ZN(G409));
  NAND3_X1  g1043(.A1(new_n994), .A2(new_n1020), .A3(G390), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G390), .B1(new_n994), .B2(new_n1020), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(new_n802), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(G390), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(G387), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT125), .B1(new_n1251), .B2(new_n1244), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1248), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1245), .B1(KEYINPUT124), .B2(new_n1246), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1246), .A2(KEYINPUT124), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1184), .A2(G378), .A3(new_n1211), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1167), .A2(new_n1170), .A3(new_n978), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1236), .B1(new_n1260), .B2(new_n1210), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1214), .A2(KEYINPUT60), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1213), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n730), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1269), .A2(KEYINPUT120), .A3(new_n1270), .A4(new_n1234), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT120), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G384), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(KEYINPUT120), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1267), .B1(new_n1214), .B2(KEYINPUT60), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1273), .B(new_n1274), .C1(new_n1275), .C2(new_n1233), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1262), .A2(new_n1263), .A3(new_n1240), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1277), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1241), .B(new_n1280), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1282));
  OAI211_X1 g1082(.A(new_n1278), .B(new_n1279), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1271), .A2(new_n1276), .A3(G2897), .A4(new_n1241), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT122), .ZN(new_n1285));
  INV_X1    g1085(.A(G2897), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1240), .B1(KEYINPUT121), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(KEYINPUT121), .B2(new_n1286), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1277), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  AOI211_X1 g1090(.A(KEYINPUT122), .B(new_n1290), .C1(new_n1271), .C2(new_n1276), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1284), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT123), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1284), .B(KEYINPUT123), .C1(new_n1289), .C2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1262), .A2(new_n1240), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1258), .B1(new_n1283), .B2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1258), .A2(KEYINPUT61), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1296), .A3(new_n1295), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1281), .A2(KEYINPUT63), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1296), .B2(new_n1280), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(G405));
  INV_X1    g1105(.A(new_n1259), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G378), .B1(new_n1184), .B2(new_n1211), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1259), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1311), .A3(new_n1277), .ZN(new_n1312));
  OAI211_X1 g1112(.A(KEYINPUT127), .B(new_n1280), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1258), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1312), .A2(new_n1258), .A3(new_n1313), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


