

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X2 U326 ( .A(n313), .B(n312), .ZN(n578) );
  XOR2_X1 U327 ( .A(n339), .B(KEYINPUT77), .Z(n294) );
  XOR2_X1 U328 ( .A(G85GAT), .B(KEYINPUT73), .Z(n295) );
  NOR2_X1 U329 ( .A1(n573), .A2(n556), .ZN(n502) );
  NOR2_X1 U330 ( .A1(n511), .A2(n510), .ZN(n512) );
  NOR2_X1 U331 ( .A1(n549), .A2(n548), .ZN(n572) );
  NOR2_X1 U332 ( .A1(n573), .A2(n566), .ZN(n554) );
  XOR2_X1 U333 ( .A(KEYINPUT28), .B(n550), .Z(n517) );
  XOR2_X1 U334 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n454) );
  XOR2_X1 U335 ( .A(KEYINPUT71), .B(KEYINPUT78), .Z(n297) );
  XNOR2_X1 U336 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n296) );
  XOR2_X1 U337 ( .A(n297), .B(n296), .Z(n313) );
  XOR2_X1 U338 ( .A(G78GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n401) );
  XOR2_X1 U341 ( .A(G64GAT), .B(KEYINPUT76), .Z(n301) );
  XNOR2_X1 U342 ( .A(G176GAT), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n435) );
  XNOR2_X1 U344 ( .A(n401), .B(n435), .ZN(n311) );
  XNOR2_X1 U345 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n302), .B(KEYINPUT75), .ZN(n303) );
  XOR2_X1 U347 ( .A(n303), .B(KEYINPUT31), .Z(n309) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G92GAT), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n295), .B(n304), .ZN(n339) );
  NAND2_X1 U350 ( .A1(G230GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n294), .B(n305), .ZN(n307) );
  XNOR2_X1 U352 ( .A(G71GAT), .B(G57GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n306), .B(KEYINPUT13), .ZN(n354) );
  XNOR2_X1 U354 ( .A(n307), .B(n354), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U357 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n315) );
  XNOR2_X1 U358 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U360 ( .A(G36GAT), .B(G50GAT), .Z(n317) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G1GAT), .Z(n415) );
  XNOR2_X1 U362 ( .A(n415), .B(KEYINPUT70), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U364 ( .A(n319), .B(n318), .Z(n321) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U367 ( .A(G22GAT), .B(G141GAT), .Z(n323) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G15GAT), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U370 ( .A(n325), .B(n324), .Z(n333) );
  XOR2_X1 U371 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n327) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(G29GAT), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U374 ( .A(KEYINPUT8), .B(n328), .Z(n348) );
  XOR2_X1 U375 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n330) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U378 ( .A(n348), .B(n331), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n573) );
  INV_X1 U380 ( .A(n573), .ZN(n532) );
  AND2_X1 U381 ( .A1(n578), .A2(n532), .ZN(n334) );
  XNOR2_X1 U382 ( .A(n334), .B(KEYINPUT79), .ZN(n466) );
  XOR2_X1 U383 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n336) );
  XNOR2_X1 U384 ( .A(KEYINPUT10), .B(KEYINPUT82), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n347) );
  XOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .Z(n432) );
  XOR2_X1 U387 ( .A(KEYINPUT9), .B(n432), .Z(n338) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(n400), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U391 ( .A(n339), .B(KEYINPUT80), .Z(n341) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U394 ( .A(n343), .B(n342), .Z(n345) );
  XNOR2_X1 U395 ( .A(G134GAT), .B(G106GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n350) );
  INV_X1 U398 ( .A(n348), .ZN(n349) );
  XOR2_X1 U399 ( .A(n350), .B(n349), .Z(n541) );
  INV_X1 U400 ( .A(n541), .ZN(n567) );
  XOR2_X1 U401 ( .A(KEYINPUT12), .B(KEYINPUT85), .Z(n356) );
  XOR2_X1 U402 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n352) );
  XNOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT83), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U407 ( .A(G8GAT), .B(G183GAT), .Z(n431) );
  XOR2_X1 U408 ( .A(G22GAT), .B(G155GAT), .Z(n399) );
  XOR2_X1 U409 ( .A(n431), .B(n399), .Z(n358) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U412 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G127GAT), .Z(n374) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U415 ( .A(G1GAT), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n374), .B(n363), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n581) );
  INV_X1 U419 ( .A(n581), .ZN(n538) );
  NAND2_X1 U420 ( .A1(n567), .A2(n538), .ZN(n368) );
  XNOR2_X1 U421 ( .A(KEYINPUT16), .B(KEYINPUT87), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n366), .B(KEYINPUT86), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n452) );
  XOR2_X1 U424 ( .A(KEYINPUT88), .B(G183GAT), .Z(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n387) );
  XOR2_X1 U427 ( .A(G176GAT), .B(G190GAT), .Z(n372) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G99GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U430 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U431 ( .A1(G227GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U433 ( .A(G71GAT), .B(KEYINPUT20), .Z(n378) );
  XNOR2_X1 U434 ( .A(G113GAT), .B(KEYINPUT89), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n385) );
  XNOR2_X1 U437 ( .A(G134GAT), .B(G120GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n381), .B(KEYINPUT0), .ZN(n424) );
  XOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n383) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n438) );
  XOR2_X1 U442 ( .A(n424), .B(n438), .Z(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U444 ( .A(n387), .B(n386), .Z(n515) );
  INV_X1 U445 ( .A(n515), .ZN(n552) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(KEYINPUT93), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(G197GAT), .B(n390), .Z(n437) );
  XOR2_X1 U450 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n392) );
  XNOR2_X1 U451 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT2), .B(KEYINPUT94), .Z(n394) );
  XNOR2_X1 U454 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n416) );
  XOR2_X1 U456 ( .A(KEYINPUT23), .B(n416), .Z(n396) );
  NAND2_X1 U457 ( .A1(G228GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n437), .B(n405), .ZN(n550) );
  NOR2_X1 U464 ( .A1(n552), .A2(n550), .ZN(n406) );
  XOR2_X1 U465 ( .A(KEYINPUT26), .B(n406), .Z(n570) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G127GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U470 ( .A(G155GAT), .B(G148GAT), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U472 ( .A(n412), .B(n411), .Z(n422) );
  XOR2_X1 U473 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U474 ( .A(KEYINPUT95), .B(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n420) );
  XOR2_X1 U476 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n423), .B(KEYINPUT96), .Z(n426) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT97), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n548) );
  INV_X1 U484 ( .A(n548), .ZN(n448) );
  NAND2_X1 U485 ( .A1(n570), .A2(n448), .ZN(n443) );
  NOR2_X1 U486 ( .A1(n552), .A2(n517), .ZN(n427) );
  NOR2_X1 U487 ( .A1(n448), .A2(n427), .ZN(n441) );
  XOR2_X1 U488 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n429) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U491 ( .A(n430), .B(G92GAT), .Z(n434) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n545) );
  XNOR2_X1 U497 ( .A(n545), .B(KEYINPUT27), .ZN(n513) );
  NOR2_X1 U498 ( .A1(n441), .A2(n513), .ZN(n442) );
  NAND2_X1 U499 ( .A1(n443), .A2(n442), .ZN(n451) );
  NOR2_X1 U500 ( .A1(n515), .A2(n545), .ZN(n444) );
  XOR2_X1 U501 ( .A(KEYINPUT100), .B(n444), .Z(n445) );
  NAND2_X1 U502 ( .A1(n550), .A2(n445), .ZN(n446) );
  XOR2_X1 U503 ( .A(KEYINPUT101), .B(n446), .Z(n447) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n447), .ZN(n449) );
  NAND2_X1 U505 ( .A1(n449), .A2(n448), .ZN(n450) );
  NAND2_X1 U506 ( .A1(n451), .A2(n450), .ZN(n461) );
  NAND2_X1 U507 ( .A1(n452), .A2(n461), .ZN(n479) );
  NOR2_X1 U508 ( .A1(n466), .A2(n479), .ZN(n459) );
  NAND2_X1 U509 ( .A1(n459), .A2(n548), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U511 ( .A(G1GAT), .B(n455), .Z(G1324GAT) );
  INV_X1 U512 ( .A(n545), .ZN(n494) );
  NAND2_X1 U513 ( .A1(n494), .A2(n459), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U515 ( .A(G15GAT), .B(KEYINPUT35), .Z(n458) );
  NAND2_X1 U516 ( .A1(n459), .A2(n552), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(G1326GAT) );
  NAND2_X1 U518 ( .A1(n517), .A2(n459), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U520 ( .A(G29GAT), .B(KEYINPUT39), .Z(n469) );
  XNOR2_X1 U521 ( .A(KEYINPUT36), .B(n567), .ZN(n585) );
  NAND2_X1 U522 ( .A1(n581), .A2(n461), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT103), .B(n462), .Z(n463) );
  NOR2_X1 U524 ( .A1(n585), .A2(n463), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT104), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT37), .ZN(n492) );
  NOR2_X1 U527 ( .A1(n492), .A2(n466), .ZN(n467) );
  XNOR2_X1 U528 ( .A(KEYINPUT38), .B(n467), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n548), .A2(n475), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(G1328GAT) );
  XOR2_X1 U531 ( .A(G36GAT), .B(KEYINPUT105), .Z(n471) );
  NAND2_X1 U532 ( .A1(n475), .A2(n494), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(G1329GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n473) );
  NAND2_X1 U535 ( .A1(n475), .A2(n552), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U537 ( .A(G43GAT), .B(n474), .Z(G1330GAT) );
  NAND2_X1 U538 ( .A1(n475), .A2(n517), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n477), .B(n578), .ZN(n534) );
  INV_X1 U543 ( .A(n534), .ZN(n556) );
  NOR2_X1 U544 ( .A1(n532), .A2(n556), .ZN(n478) );
  XOR2_X1 U545 ( .A(KEYINPUT108), .B(n478), .Z(n491) );
  NOR2_X1 U546 ( .A1(n491), .A2(n479), .ZN(n480) );
  XOR2_X1 U547 ( .A(KEYINPUT109), .B(n480), .Z(n487) );
  NAND2_X1 U548 ( .A1(n487), .A2(n548), .ZN(n481) );
  XNOR2_X1 U549 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U550 ( .A(G57GAT), .B(n483), .ZN(G1332GAT) );
  NAND2_X1 U551 ( .A1(n494), .A2(n487), .ZN(n484) );
  XNOR2_X1 U552 ( .A(n484), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U553 ( .A1(n552), .A2(n487), .ZN(n485) );
  XNOR2_X1 U554 ( .A(n485), .B(KEYINPUT110), .ZN(n486) );
  XNOR2_X1 U555 ( .A(G71GAT), .B(n486), .ZN(G1334GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n489) );
  NAND2_X1 U557 ( .A1(n487), .A2(n517), .ZN(n488) );
  XNOR2_X1 U558 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U559 ( .A(G78GAT), .B(n490), .Z(G1335GAT) );
  NOR2_X1 U560 ( .A1(n492), .A2(n491), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n499), .A2(n548), .ZN(n493) );
  XNOR2_X1 U562 ( .A(n493), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U563 ( .A1(n494), .A2(n499), .ZN(n495) );
  XNOR2_X1 U564 ( .A(n495), .B(KEYINPUT112), .ZN(n496) );
  XNOR2_X1 U565 ( .A(G92GAT), .B(n496), .ZN(G1337GAT) );
  XOR2_X1 U566 ( .A(G99GAT), .B(KEYINPUT113), .Z(n498) );
  NAND2_X1 U567 ( .A1(n499), .A2(n552), .ZN(n497) );
  XNOR2_X1 U568 ( .A(n498), .B(n497), .ZN(G1338GAT) );
  NAND2_X1 U569 ( .A1(n517), .A2(n499), .ZN(n500) );
  XNOR2_X1 U570 ( .A(n500), .B(KEYINPUT44), .ZN(n501) );
  XNOR2_X1 U571 ( .A(G106GAT), .B(n501), .ZN(G1339GAT) );
  XOR2_X1 U572 ( .A(n581), .B(KEYINPUT114), .Z(n561) );
  XNOR2_X1 U573 ( .A(n502), .B(KEYINPUT46), .ZN(n503) );
  NOR2_X1 U574 ( .A1(n561), .A2(n503), .ZN(n504) );
  NAND2_X1 U575 ( .A1(n504), .A2(n567), .ZN(n505) );
  XNOR2_X1 U576 ( .A(KEYINPUT47), .B(n505), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n507) );
  NOR2_X1 U578 ( .A1(n585), .A2(n581), .ZN(n506) );
  XNOR2_X1 U579 ( .A(n507), .B(n506), .ZN(n509) );
  NAND2_X1 U580 ( .A1(n578), .A2(n573), .ZN(n508) );
  NOR2_X1 U581 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U582 ( .A(KEYINPUT48), .B(n512), .ZN(n544) );
  NOR2_X1 U583 ( .A1(n544), .A2(n513), .ZN(n514) );
  NAND2_X1 U584 ( .A1(n548), .A2(n514), .ZN(n530) );
  NOR2_X1 U585 ( .A1(n515), .A2(n530), .ZN(n516) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(n516), .Z(n518) );
  NOR2_X1 U587 ( .A1(n518), .A2(n517), .ZN(n523) );
  INV_X1 U588 ( .A(n523), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n573), .A2(n526), .ZN(n520) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n519) );
  XNOR2_X1 U591 ( .A(n520), .B(n519), .ZN(G1340GAT) );
  NOR2_X1 U592 ( .A1(n556), .A2(n526), .ZN(n522) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n521) );
  XNOR2_X1 U594 ( .A(n522), .B(n521), .ZN(G1341GAT) );
  NAND2_X1 U595 ( .A1(n523), .A2(n561), .ZN(n524) );
  XNOR2_X1 U596 ( .A(n524), .B(KEYINPUT50), .ZN(n525) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n525), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n567), .A2(n526), .ZN(n528) );
  XNOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n529), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n570), .A2(n530), .ZN(n531) );
  XOR2_X1 U603 ( .A(KEYINPUT119), .B(n531), .Z(n540) );
  NAND2_X1 U604 ( .A1(n540), .A2(n532), .ZN(n533) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n533), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n536) );
  NAND2_X1 U607 ( .A1(n540), .A2(n534), .ZN(n535) );
  XNOR2_X1 U608 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(n537), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n540), .A2(n538), .ZN(n539) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(n539), .ZN(G1346GAT) );
  XNOR2_X1 U612 ( .A(G162GAT), .B(KEYINPUT120), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U614 ( .A(n543), .B(n542), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U616 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n546) );
  XNOR2_X1 U617 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n572), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT55), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n566) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n555), .ZN(G1348GAT) );
  NOR2_X1 U623 ( .A1(n566), .A2(n556), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  INV_X1 U628 ( .A(n566), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n565) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(n569), .B(n568), .Z(G1351GAT) );
  INV_X1 U636 ( .A(n570), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n584) );
  NOR2_X1 U638 ( .A1(n573), .A2(n584), .ZN(n577) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n584), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

