//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT68), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n479), .A2(G137), .A3(new_n465), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND3_X1  g058(.A1(new_n479), .A2(G2105), .A3(new_n480), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n480), .A2(new_n478), .A3(new_n465), .A4(new_n469), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n480), .A2(new_n478), .A3(new_n469), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n467), .A2(new_n469), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n480), .A2(new_n478), .A3(new_n469), .A4(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n506), .B2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT72), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(KEYINPUT73), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n514), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n516), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT6), .A3(new_n510), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n520), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND4_X1   g104(.A1(new_n525), .A2(new_n518), .A3(new_n529), .A4(new_n517), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n511), .A2(new_n512), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n529), .A2(G62), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT74), .Z(new_n536));
  OAI21_X1  g111(.A(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n522), .A2(new_n531), .A3(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND2_X1  g114(.A1(new_n521), .A2(G51), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(G89), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AND2_X1   g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n529), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(new_n521), .A2(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n532), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n530), .A2(G90), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n521), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n532), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n530), .A2(G81), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g136(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n521), .A2(new_n566), .A3(G53), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n525), .A2(G543), .A3(new_n518), .A4(new_n517), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g146(.A1(KEYINPUT76), .A2(G65), .ZN(new_n572));
  NAND2_X1  g147(.A1(KEYINPUT76), .A2(G65), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n529), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n516), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G91), .B2(new_n530), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  AND2_X1   g154(.A1(new_n527), .A2(new_n528), .ZN(new_n580));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n516), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n521), .B2(G49), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT77), .B1(new_n530), .B2(G87), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n525), .A2(new_n529), .A3(new_n518), .A4(new_n517), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n583), .B1(new_n584), .B2(new_n588), .ZN(G288));
  NOR2_X1   g164(.A1(new_n514), .A2(new_n519), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n590), .A2(G86), .A3(new_n529), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n527), .B2(new_n528), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n533), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n517), .A2(new_n518), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n596), .A2(G48), .A3(G543), .A4(new_n525), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n595), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n532), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT78), .Z(new_n601));
  AOI22_X1  g176(.A1(G47), .A2(new_n521), .B1(new_n530), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n585), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n516), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n568), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n558), .A2(new_n619), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n615), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n619), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n492), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n465), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n633), .C2(new_n484), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n498), .A2(new_n473), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n636), .A2(G2096), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n640), .B1(new_n644), .B2(G2100), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n637), .A2(new_n642), .A3(new_n643), .A4(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n667), .A2(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(KEYINPUT85), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(new_n673), .A3(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n667), .B(KEYINPUT17), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n665), .C1(new_n675), .C2(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n669), .A3(new_n664), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n671), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(KEYINPUT87), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  NOR3_X1   g266(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  XNOR2_X1  g277(.A(KEYINPUT31), .B(G11), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT30), .B(G28), .Z(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NOR2_X1   g280(.A1(G171), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G5), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n703), .B1(G29), .B2(new_n704), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G168), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G16), .B2(G21), .ZN(new_n711));
  INV_X1    g286(.A(G1966), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n636), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n709), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT96), .Z(new_n718));
  AND2_X1   g293(.A1(new_n715), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n492), .A2(G141), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n724), .A2(new_n725), .B1(G105), .B2(new_n473), .ZN(new_n726));
  INV_X1    g301(.A(G129), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n484), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n721), .A2(KEYINPUT94), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n719), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT95), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n718), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G162), .A2(G29), .ZN(new_n740));
  OR2_X1    g315(.A1(G29), .A2(G35), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n715), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n492), .A2(G140), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(new_n484), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G128), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n715), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n498), .A2(G127), .ZN(new_n760));
  INV_X1    g335(.A(G115), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n466), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  NAND2_X1  g338(.A1(G103), .A2(G2104), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n762), .A2(G2105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n492), .A2(G139), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n759), .B1(new_n769), .B2(new_n715), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n482), .B2(new_n715), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n770), .A2(G2072), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G2072), .B2(new_n770), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n705), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n705), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n559), .B2(new_n705), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n777), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n745), .A2(new_n758), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n707), .A2(new_n708), .B1(new_n771), .B2(new_n775), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n735), .B2(new_n736), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT97), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n705), .A2(G4), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n616), .B2(new_n705), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1348), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n715), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n715), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n792), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n739), .A2(new_n786), .A3(new_n789), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n705), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n705), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT90), .Z(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n804), .A2(new_n805), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G23), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT89), .Z(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G288), .B2(new_n705), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n806), .A2(new_n809), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n705), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n705), .B2(G24), .ZN(new_n821));
  INV_X1    g396(.A(G1986), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n715), .A2(G25), .ZN(new_n825));
  INV_X1    g400(.A(G119), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n465), .A2(G107), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n484), .A2(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n492), .A2(G131), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n715), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT88), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n823), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n817), .A2(new_n818), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n838));
  OR2_X1    g413(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n838), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n801), .A2(new_n840), .A3(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  NAND2_X1  g418(.A1(new_n521), .A2(G55), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n530), .A2(G93), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n844), .B(new_n845), .C1(new_n532), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n616), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n559), .B(new_n847), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(KEYINPUT38), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n847), .B(new_n558), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT100), .Z(new_n859));
  AOI21_X1  g434(.A(KEYINPUT39), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n849), .B1(new_n859), .B2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(KEYINPUT105), .B(G37), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n769), .A2(KEYINPUT102), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT101), .Z(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n734), .A2(new_n755), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n498), .A2(new_n499), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n505), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n755), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n732), .A2(new_n733), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n868), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n867), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n866), .A3(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n492), .A2(G142), .ZN(new_n885));
  OR2_X1    g460(.A1(G106), .A2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n887));
  INV_X1    g462(.A(G130), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n885), .B(new_n887), .C1(new_n888), .C2(new_n484), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n639), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n639), .A2(new_n889), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(new_n831), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n831), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n636), .B(new_n482), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(G162), .Z(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n884), .B2(new_n894), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n864), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n884), .A2(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n884), .A2(new_n897), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n884), .A2(new_n906), .A3(new_n897), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n900), .ZN(new_n909));
  OAI211_X1 g484(.A(KEYINPUT40), .B(new_n902), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n884), .A2(new_n906), .A3(new_n897), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n906), .B1(new_n884), .B2(new_n897), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n898), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n900), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n915), .B2(new_n902), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n911), .A2(new_n916), .ZN(G395));
  NAND2_X1  g492(.A1(new_n847), .A2(new_n619), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  XNOR2_X1  g494(.A(G288), .B(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G290), .ZN(new_n921));
  XOR2_X1   g496(.A(G303), .B(G305), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  INV_X1    g502(.A(G299), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n615), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n615), .A2(KEYINPUT107), .A3(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT108), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n856), .B(KEYINPUT106), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(new_n626), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n926), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n918), .B1(new_n943), .B2(new_n619), .ZN(G295));
  OAI21_X1  g519(.A(new_n918), .B1(new_n943), .B2(new_n619), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n853), .A2(G301), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n856), .A2(G171), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n947), .A2(new_n948), .A3(G286), .ZN(new_n949));
  OAI21_X1  g524(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n938), .A2(new_n940), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(G303), .B(G305), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n921), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n937), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n923), .A2(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n959), .A2(new_n961), .B1(new_n951), .B2(new_n955), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n946), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n933), .A2(new_n954), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n951), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n863), .A3(new_n956), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n968), .B2(new_n946), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT44), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n967), .A2(new_n946), .A3(new_n863), .A4(new_n956), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT43), .B1(new_n958), .B2(new_n962), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(KEYINPUT118), .ZN(new_n977));
  NOR2_X1   g552(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(G164), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n470), .A2(new_n471), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G2105), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n481), .A2(new_n982), .A3(G40), .A4(new_n474), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n500), .B2(new_n505), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n507), .B1(new_n502), .B2(new_n504), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n871), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT118), .A3(new_n978), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n980), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1956), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT112), .B(G1384), .Z(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n871), .B2(new_n872), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n983), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1002), .B(new_n1003), .C1(new_n571), .C2(new_n577), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n571), .A2(new_n577), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1001), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n985), .A2(new_n983), .A3(G2067), .ZN(new_n1011));
  INV_X1    g586(.A(G137), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n491), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G40), .ZN(new_n1014));
  NOR4_X1   g589(.A1(new_n1013), .A2(new_n472), .A3(new_n1014), .A4(new_n475), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n984), .C1(new_n500), .C2(new_n505), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n506), .A2(new_n508), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n1018), .B2(new_n871), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1015), .B(new_n1017), .C1(new_n1019), .C2(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(G1348), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1011), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT121), .B1(new_n1022), .B2(new_n615), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1017), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n989), .A2(new_n984), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1348), .B1(new_n1027), .B2(new_n1015), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1024), .B(new_n616), .C1(new_n1028), .C2(new_n1011), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1010), .A2(new_n1023), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1008), .A2(new_n993), .A3(new_n1000), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT61), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1008), .A2(new_n993), .A3(new_n1000), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1008), .B1(new_n993), .B2(new_n1000), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n1031), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT58), .B(G1341), .Z(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n985), .B2(new_n983), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT122), .B(new_n1039), .C1(new_n985), .C2(new_n983), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n989), .B2(new_n984), .ZN(new_n1045));
  INV_X1    g620(.A(new_n996), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT45), .B(new_n1046), .C1(new_n500), .C2(new_n505), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1015), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1045), .A2(new_n1048), .A3(G1996), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n559), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g628(.A(new_n559), .B1(KEYINPUT123), .B2(new_n1051), .C1(new_n1044), .C2(new_n1049), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1028), .B2(new_n1011), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1022), .A2(KEYINPUT60), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n616), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1022), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1032), .B1(new_n1038), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n995), .A2(new_n998), .A3(new_n795), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT124), .B(G1961), .Z(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1065), .B1(new_n1020), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(G164), .A2(new_n994), .A3(G1384), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1384), .B1(new_n871), .B2(new_n872), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1015), .B1(new_n1069), .B2(KEYINPUT45), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n795), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1065), .A2(new_n1064), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1020), .A2(new_n1066), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1064), .B(G2078), .C1(new_n983), .C2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n997), .A2(KEYINPUT45), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1015), .A2(KEYINPUT125), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1047), .A4(new_n1079), .ZN(new_n1080));
  AND4_X1   g655(.A1(G301), .A2(new_n1074), .A3(new_n1075), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1063), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1074), .A2(new_n1075), .A3(new_n1080), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1067), .A2(G301), .A3(new_n1072), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(KEYINPUT54), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n712), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n983), .A2(G2084), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1017), .B(new_n1088), .C1(new_n1019), .C2(new_n1016), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1089), .A3(G168), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1090), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1082), .A2(new_n1086), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G303), .A2(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1016), .B1(new_n989), .B2(new_n984), .ZN(new_n1104));
  NOR4_X1   g679(.A1(new_n1104), .A2(new_n1025), .A3(G2090), .A4(new_n983), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1971), .B1(new_n995), .B2(new_n998), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1069), .B2(new_n1015), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT115), .B(G86), .Z(new_n1110));
  NAND4_X1  g685(.A1(new_n596), .A2(new_n525), .A3(new_n529), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n597), .A2(new_n1111), .A3(new_n595), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G1981), .ZN(new_n1113));
  INV_X1    g688(.A(G1981), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n591), .A2(new_n597), .A3(new_n1114), .A4(new_n595), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1115), .A3(KEYINPUT116), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT49), .B1(new_n1116), .B2(KEYINPUT117), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(KEYINPUT117), .B2(KEYINPUT49), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1109), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1976), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G288), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n590), .A2(KEYINPUT77), .A3(G87), .A4(new_n529), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(G1976), .A3(new_n583), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1123), .A2(new_n1109), .A3(new_n1124), .A4(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1127), .A2(G1976), .A3(new_n583), .ZN(new_n1130));
  OAI21_X1  g705(.A(G8), .B1(new_n985), .B2(new_n983), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT52), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1107), .A2(new_n1121), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G2090), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n980), .A2(new_n986), .A3(new_n1135), .A4(new_n990), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n805), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1103), .B1(new_n1138), .B2(G8), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1098), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT49), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1120), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1146), .B2(new_n1109), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(G8), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1103), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT126), .A4(new_n1107), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1140), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1062), .A2(new_n1097), .A3(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1108), .B(G286), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1147), .A2(new_n1150), .A3(new_n1107), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1107), .A2(new_n1121), .A3(new_n1133), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1158), .A2(KEYINPUT119), .A3(new_n1150), .A4(new_n1154), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(G8), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1149), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1158), .A2(KEYINPUT63), .A3(new_n1154), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1073), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1096), .B2(KEYINPUT62), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1152), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1107), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1127), .A2(new_n1122), .A3(new_n583), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1115), .B1(new_n1146), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1170), .A2(new_n1147), .B1(new_n1172), .B2(new_n1109), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1153), .A2(new_n1165), .A3(new_n1169), .A4(new_n1173), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1078), .A2(KEYINPUT113), .A3(new_n983), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT113), .B1(new_n1078), .B2(new_n983), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n734), .A2(G1996), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n1177), .A2(new_n1178), .A3(KEYINPUT114), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT114), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1177), .ZN(new_n1182));
  INV_X1    g757(.A(new_n831), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1183), .A2(new_n834), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n834), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n734), .A2(G1996), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n755), .B(G2067), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1181), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n819), .A2(new_n822), .ZN(new_n1191));
  NAND2_X1  g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1177), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1174), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1177), .A2(new_n1196), .A3(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1182), .B1(new_n734), .B2(new_n1188), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1196), .B1(new_n1177), .B2(G1996), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(KEYINPUT47), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(KEYINPUT47), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  OAI22_X1  g779(.A1(new_n1201), .A2(new_n1202), .B1(new_n1190), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1181), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n874), .A2(new_n757), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1177), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1195), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1195), .A2(KEYINPUT127), .A3(new_n1209), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g789(.A(new_n662), .ZN(new_n1216));
  NOR3_X1   g790(.A1(new_n1216), .A2(new_n463), .A3(G227), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n701), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n1218), .B1(new_n971), .B2(new_n972), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n915), .A2(new_n902), .ZN(new_n1220));
  AND2_X1   g794(.A1(new_n1219), .A2(new_n1220), .ZN(G308));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(G225));
endmodule


