//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G234));
  NAND2_X1  g028(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  AOI22_X1  g037(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n473), .A2(KEYINPUT70), .A3(G137), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n469), .A2(KEYINPUT71), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n470), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(KEYINPUT72), .A3(G124), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n484), .A2(new_n486), .A3(new_n470), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n491), .A2(new_n492), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(G102), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n476), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n466), .A3(new_n468), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n473), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(G543), .A3(new_n523), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n522), .A2(G62), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT74), .ZN(new_n532));
  OAI21_X1  g107(.A(G651), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n529), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n525), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI211_X1 g117(.A(new_n540), .B(new_n541), .C1(new_n522), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n515), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n525), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n528), .A2(G52), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(G81), .A2(new_n525), .B1(new_n528), .B2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n521), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G651), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n527), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n527), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n525), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n521), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(G299));
  OR2_X1    g151(.A1(G171), .A2(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(G171), .A2(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G301));
  NAND2_X1  g154(.A1(new_n525), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n528), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n521), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n527), .B2(new_n588), .C1(new_n589), .C2(new_n524), .ZN(G305));
  NAND2_X1  g165(.A1(new_n525), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n528), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n515), .C2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n578), .B2(new_n577), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n525), .A2(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G79), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT79), .B1(new_n600), .B2(new_n518), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n600), .A2(new_n518), .A3(KEYINPUT79), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n521), .C2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n596), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT78), .B2(new_n596), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(KEYINPUT78), .B2(new_n596), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n611), .B1(new_n613), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n606), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n559), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n619), .B(new_n620), .S(KEYINPUT81), .Z(G323));
  XOR2_X1   g196(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  NAND2_X1  g198(.A1(new_n473), .A2(new_n477), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2100), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n488), .A2(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n494), .A2(G135), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n660), .A2(KEYINPUT17), .A3(new_n657), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n660), .B2(KEYINPUT17), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n661), .A2(new_n662), .A3(new_n656), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT85), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n667), .A2(new_n668), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n672), .A3(new_n675), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G4), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n606), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1348), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(G21), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G168), .B2(new_n690), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT94), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G1966), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n494), .A2(G139), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n477), .A2(G103), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT25), .Z(new_n700));
  AOI22_X1  g275(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n700), .C1(new_n470), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G33), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G2072), .Z(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  AND2_X1   g280(.A1(KEYINPUT24), .A2(G34), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(KEYINPUT24), .B2(G34), .ZN(new_n707));
  OAI22_X1  g282(.A1(G160), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G2084), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n632), .A2(new_n705), .ZN(new_n710));
  INV_X1    g285(.A(G28), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n713));
  OR2_X1    g288(.A1(KEYINPUT31), .A2(G11), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n704), .A2(new_n709), .A3(new_n710), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G171), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G5), .B2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n488), .A2(G129), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n494), .A2(G141), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT26), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n477), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  OAI22_X1  g307(.A1(new_n719), .A2(new_n720), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OR4_X1    g308(.A1(new_n693), .A2(new_n697), .A3(new_n717), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G164), .A2(new_n705), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n705), .A2(G27), .ZN(new_n736));
  OAI21_X1  g311(.A(KEYINPUT96), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT96), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT97), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n719), .A2(new_n720), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G2084), .B2(new_n708), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n731), .B2(new_n732), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT95), .Z(new_n745));
  NOR3_X1   g320(.A1(new_n734), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n705), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n705), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n690), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n559), .B2(new_n690), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n690), .A2(G20), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n756), .B(new_n757), .C1(G299), .C2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  INV_X1    g334(.A(G1956), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n751), .A2(new_n755), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n488), .A2(G128), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G140), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n493), .A2(KEYINPUT92), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT92), .B1(new_n493), .B2(new_n767), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n766), .A2(KEYINPUT93), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n768), .A2(new_n763), .A3(new_n769), .A4(new_n765), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n705), .ZN(new_n776));
  INV_X1    g351(.A(G26), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT28), .B2(new_n778), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n762), .B1(G2067), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n746), .B(new_n781), .C1(G2067), .C2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n690), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n690), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n690), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n690), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G6), .B(G305), .S(G16), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n786), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT34), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n705), .A2(G25), .ZN(new_n798));
  INV_X1    g373(.A(G131), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n493), .A2(KEYINPUT89), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n488), .A2(G119), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT89), .B1(new_n493), .B2(new_n799), .ZN(new_n802));
  OR2_X1    g377(.A1(G95), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n798), .B1(new_n806), .B2(new_n705), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1986), .Z(new_n812));
  NAND3_X1  g387(.A1(new_n797), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT36), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n782), .A2(new_n814), .ZN(G311));
  INV_X1    g390(.A(G311), .ZN(G150));
  NAND2_X1  g391(.A1(new_n606), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n525), .A2(G93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n528), .A2(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n820), .B(new_n821), .C1(new_n515), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n559), .B(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n819), .A2(new_n824), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n825), .A2(new_n826), .A3(G860), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(G860), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  NAND3_X1  g405(.A1(new_n770), .A2(new_n806), .A3(new_n773), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n806), .B1(new_n770), .B2(new_n773), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n625), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n833), .ZN(new_n835));
  INV_X1    g410(.A(new_n625), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n831), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n488), .A2(G130), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n494), .A2(G142), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n840), .A2(new_n470), .A3(G118), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n470), .B2(G118), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n838), .B(new_n839), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n702), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n834), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n834), .B2(new_n837), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n505), .A2(new_n849), .A3(new_n512), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n505), .B2(new_n512), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n834), .A2(new_n837), .ZN(new_n855));
  INV_X1    g430(.A(new_n845), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n854), .B1(new_n857), .B2(new_n846), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n729), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n852), .B1(new_n847), .B2(new_n848), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n854), .A3(new_n846), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n730), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT102), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n859), .B2(new_n862), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n498), .B(G160), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n632), .B(KEYINPUT98), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OAI22_X1  g443(.A1(KEYINPUT101), .A2(new_n863), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n859), .A2(new_n862), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n864), .B(new_n870), .C1(new_n871), .C2(KEYINPUT102), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT40), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n869), .A2(new_n872), .A3(new_n876), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(G395));
  OR2_X1    g453(.A1(new_n618), .A2(new_n824), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n618), .A2(new_n824), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n612), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n606), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n612), .A2(new_n883), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n606), .A2(new_n883), .A3(new_n612), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n606), .A3(new_n884), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n881), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n879), .A2(new_n880), .A3(new_n890), .A4(new_n892), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n788), .B(G290), .ZN(new_n902));
  XOR2_X1   g477(.A(G303), .B(G305), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n899), .B2(KEYINPUT42), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT42), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n901), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n823), .A2(new_n595), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(G331));
  INV_X1    g487(.A(new_n824), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(G168), .ZN(new_n914));
  NAND2_X1  g489(.A1(G171), .A2(G286), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n915), .B(KEYINPUT106), .ZN(new_n919));
  AOI21_X1  g494(.A(G286), .B1(new_n577), .B2(new_n578), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n824), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n893), .A3(new_n889), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n918), .A2(new_n921), .A3(new_n890), .A4(new_n892), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n904), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  INV_X1    g503(.A(new_n904), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n904), .A4(new_n924), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n930), .A3(new_n873), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT109), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n927), .A2(new_n873), .A3(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n904), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n937), .B2(new_n928), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(KEYINPUT44), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n933), .A2(KEYINPUT109), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n935), .B2(new_n939), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n941), .A2(new_n942), .B1(new_n945), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g521(.A(new_n503), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n473), .B2(G126), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n948), .A2(new_n470), .B1(new_n500), .B2(new_n476), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n510), .B1(new_n473), .B2(new_n507), .ZN(new_n950));
  AND4_X1   g525(.A1(new_n510), .A2(new_n507), .A3(new_n466), .A4(new_n468), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT99), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n505), .A2(new_n849), .A3(new_n512), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n479), .A2(G40), .A3(new_n481), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n774), .B(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n729), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT112), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n805), .A2(new_n808), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n775), .A2(new_n962), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n960), .A2(new_n964), .ZN(new_n972));
  NAND2_X1  g547(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n972), .B(new_n973), .Z(new_n974));
  AND2_X1   g549(.A1(new_n963), .A2(new_n730), .ZN(new_n975));
  OAI221_X1 g550(.A(new_n974), .B1(KEYINPUT127), .B2(KEYINPUT46), .C1(new_n975), .C2(new_n961), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  NOR2_X1   g552(.A1(new_n806), .A2(new_n809), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n960), .B1(new_n968), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT110), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n960), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n971), .B(new_n977), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g561(.A1(G286), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT123), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n986), .B(KEYINPUT51), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AND4_X1   g564(.A1(G40), .A2(new_n481), .A3(new_n478), .A4(new_n475), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n949), .B2(new_n952), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n957), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n513), .B2(new_n991), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT115), .B(G1384), .C1(new_n505), .C2(new_n512), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n993), .B1(new_n957), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n959), .B1(KEYINPUT50), .B2(new_n992), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(KEYINPUT50), .B2(new_n997), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n998), .A2(G1966), .B1(new_n1000), .B2(G2084), .ZN(new_n1001));
  OAI211_X1 g576(.A(G8), .B(new_n989), .C1(new_n1001), .C2(G286), .ZN(new_n1002));
  INV_X1    g577(.A(new_n987), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1001), .A2(new_n1003), .B1(new_n986), .B2(KEYINPUT51), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1001), .B2(G8), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n988), .B2(KEYINPUT51), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n992), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n505), .B2(new_n512), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1014), .A3(new_n990), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n991), .C1(new_n850), .C2(new_n851), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n955), .A2(new_n1018), .A3(KEYINPUT45), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1010), .B1(new_n1021), .B2(G2078), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1000), .A2(new_n720), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n998), .A2(KEYINPUT53), .A3(new_n740), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G301), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1009), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G305), .B(G1981), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n997), .A2(new_n959), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n788), .A2(G1976), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT55), .Z(new_n1047));
  NOR2_X1   g622(.A1(new_n1020), .A2(G1971), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1000), .A2(G2090), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1047), .B(G8), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1048), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n992), .A2(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1013), .A2(new_n994), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(KEYINPUT50), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n990), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(KEYINPUT116), .A3(new_n990), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n750), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1034), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1045), .B(new_n1050), .C1(new_n1047), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT126), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1027), .B(new_n1029), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1037), .A2(new_n1041), .A3(new_n788), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G305), .A2(G1981), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1035), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1050), .B2(new_n1044), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1001), .A2(G8), .A3(G168), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1047), .B1(new_n1074), .B2(G8), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1075), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n1050), .A3(new_n1045), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1070), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1066), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1025), .B2(G301), .ZN(new_n1081));
  INV_X1    g656(.A(G171), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n479), .A2(KEYINPUT125), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n479), .A2(KEYINPUT125), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n481), .A2(KEYINPUT53), .A3(G40), .A4(new_n740), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1018), .B1(new_n955), .B2(KEYINPUT45), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n958), .B(new_n1086), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1022), .A2(new_n1023), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1081), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1022), .A2(G301), .A3(new_n1023), .A4(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1025), .B2(G301), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1093), .A2(new_n1080), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1091), .B(new_n1094), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n612), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n995), .A2(new_n996), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1057), .B1(new_n1103), .B2(new_n959), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1052), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1059), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n760), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1109), .A3(new_n760), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT56), .B(G2072), .Z(new_n1112));
  NOR2_X1   g687(.A1(new_n1021), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1101), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g690(.A(KEYINPUT117), .B(G1956), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1109), .B1(new_n1106), .B2(new_n760), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1101), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1000), .A2(new_n1119), .B1(new_n1033), .B2(new_n962), .ZN(new_n1120));
  INV_X1    g695(.A(new_n606), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1118), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(KEYINPUT60), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(new_n606), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(KEYINPUT60), .B2(new_n1120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1011), .A2(new_n1014), .A3(new_n990), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n964), .B(new_n1133), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n990), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT119), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1134), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1132), .B1(new_n1144), .B2(new_n559), .ZN(new_n1145));
  AOI211_X1 g720(.A(KEYINPUT119), .B(new_n1138), .C1(new_n1020), .C2(new_n964), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1132), .B(new_n559), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1131), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1100), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n559), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT59), .A3(new_n1148), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1150), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1123), .B1(new_n1130), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1095), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(KEYINPUT121), .B(new_n1123), .C1(new_n1130), .C2(new_n1157), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1079), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n960), .A2(G1986), .A3(G290), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n983), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT111), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n980), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n985), .B1(new_n1162), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g742(.A(G319), .ZN(new_n1169));
  NOR4_X1   g743(.A1(G401), .A2(G229), .A3(new_n1169), .A4(G227), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n1170), .B1(new_n943), .B2(new_n944), .ZN(new_n1171));
  AND2_X1   g745(.A1(new_n869), .A2(new_n873), .ZN(new_n1172));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1172), .B2(new_n872), .ZN(G308));
  OAI211_X1 g747(.A(new_n874), .B(new_n1170), .C1(new_n943), .C2(new_n944), .ZN(G225));
endmodule


