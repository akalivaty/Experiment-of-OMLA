//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT67), .B(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n202), .A2(G50), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n218), .A2(KEYINPUT1), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(new_n209), .B2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n208), .A2(KEYINPUT65), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n223), .B(new_n231), .C1(KEYINPUT1), .C2(new_n218), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XOR2_X1   g0044(.A(G58), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(new_n210), .B2(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n258), .A2(new_n272), .A3(new_n267), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n219), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n281), .A3(new_n219), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT8), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n207), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n207), .B1(new_n201), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n283), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n280), .A2(new_n298), .A3(new_n282), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n207), .A2(G1), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(G50), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n295), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n297), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n277), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n275), .A2(G200), .B1(new_n305), .B2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n275), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n305), .C1(G179), .C2(new_n275), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(new_n292), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n319), .B1(new_n207), .B2(new_n210), .C1(new_n290), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n321), .A2(new_n279), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n301), .A2(G77), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n298), .A2(new_n219), .A3(new_n278), .ZN(new_n324));
  INV_X1    g0124(.A(new_n210), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n298), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n258), .A2(new_n272), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n262), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n211), .B2(new_n269), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT72), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n333));
  INV_X1    g0133(.A(G107), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(new_n334), .B2(new_n252), .C1(new_n255), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n258), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n331), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n327), .B1(new_n339), .B2(new_n276), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n338), .A2(new_n337), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n332), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n339), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n327), .B1(new_n339), .B2(new_n315), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n318), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G68), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n324), .A2(new_n352), .A3(new_n300), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n206), .A2(new_n352), .A3(G13), .A4(G20), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT12), .B1(new_n354), .B2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(KEYINPUT74), .A3(KEYINPUT12), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n352), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n290), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n283), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT11), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n283), .A2(new_n362), .A3(KEYINPUT11), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n367), .A2(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n269), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n264), .A2(KEYINPUT73), .A3(new_n268), .A4(new_n266), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G238), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n238), .A2(G1698), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G226), .B2(G1698), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n273), .B1(new_n383), .B2(new_n258), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n375), .A2(new_n376), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n376), .B1(new_n375), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g0186(.A(G169), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(new_n376), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n387), .A2(KEYINPUT14), .B1(new_n391), .B2(new_n346), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n391), .B2(G169), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n371), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G200), .B1(new_n385), .B2(new_n386), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n370), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT76), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n399), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n288), .A2(new_n301), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n280), .A2(new_n298), .A3(new_n282), .ZN(new_n406));
  AOI221_X4 g0206(.A(KEYINPUT77), .B1(new_n405), .B2(new_n298), .C1(new_n406), .C2(new_n288), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n288), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n298), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  OR2_X1    g0213(.A1(KEYINPUT3), .A2(G33), .ZN(new_n414));
  NAND2_X1  g0214(.A1(KEYINPUT3), .A2(G33), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n207), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n415), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n352), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n284), .A2(new_n352), .ZN(new_n421));
  OAI21_X1  g0221(.A(G20), .B1(new_n421), .B2(new_n201), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n292), .A2(G159), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n413), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n382), .B2(new_n207), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n380), .A2(new_n381), .A3(new_n417), .A4(G20), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n424), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(KEYINPUT16), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n430), .A3(new_n279), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n412), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G223), .A2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n270), .B2(G1698), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n252), .B1(G33), .B2(G87), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(new_n266), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n264), .A2(G232), .A3(new_n268), .A4(new_n266), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(G190), .A3(new_n329), .A4(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n329), .B(new_n437), .C1(new_n435), .C2(new_n266), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n404), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n438), .A2(new_n440), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n431), .A4(new_n412), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(G169), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n436), .A2(G179), .A3(new_n329), .A4(new_n437), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n412), .A2(new_n431), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n446), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n425), .A2(new_n430), .A3(new_n279), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n409), .A2(new_n410), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT77), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n409), .A2(new_n408), .A3(new_n410), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n460), .B2(new_n449), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n445), .B1(new_n451), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n351), .A2(new_n400), .A3(new_n403), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(G33), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G116), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n324), .A2(new_n465), .B1(G116), .B2(new_n298), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n207), .C1(G33), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT20), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  AOI22_X1  g0271(.A1(KEYINPUT85), .A2(new_n470), .B1(new_n471), .B2(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n472), .A3(new_n279), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n469), .A2(new_n472), .A3(new_n474), .A4(new_n279), .ZN(new_n477));
  AOI211_X1 g0277(.A(KEYINPUT86), .B(new_n466), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  INV_X1    g0280(.A(new_n466), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(G169), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G264), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(new_n253), .C1(new_n380), .C2(new_n381), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n414), .A2(G303), .A3(new_n415), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n487), .A2(new_n258), .ZN(new_n488));
  OR2_X1    g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n261), .A2(G1), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(G274), .A3(new_n266), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n490), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n266), .ZN(new_n497));
  INV_X1    g0297(.A(G270), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT84), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n206), .A2(G45), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n489), .B2(new_n490), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n258), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G270), .B1(new_n328), .B2(new_n502), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n487), .A2(new_n258), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n483), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n480), .A2(new_n481), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n480), .A2(new_n479), .A3(new_n481), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n504), .A2(G179), .A3(new_n506), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n509), .A2(KEYINPUT21), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(G190), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n517), .B(new_n518), .C1(new_n341), .C2(new_n508), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT87), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n499), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n513), .A3(G169), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n520), .B(new_n525), .C1(new_n483), .C2(new_n508), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n516), .B(new_n519), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(new_n253), .C1(new_n380), .C2(new_n381), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n252), .A2(G244), .A3(new_n253), .A4(new_n532), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n467), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n258), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  INV_X1    g0339(.A(G257), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n493), .B1(new_n497), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n539), .B1(new_n538), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n315), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n546), .A2(new_n468), .A3(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(G97), .B(G107), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n549), .A2(new_n207), .B1(new_n361), .B2(new_n293), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n334), .B1(new_n418), .B2(new_n419), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n279), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n303), .A2(G97), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n280), .A2(new_n298), .A3(new_n464), .A4(new_n282), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(KEYINPUT79), .B(new_n553), .C1(new_n554), .C2(G97), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n538), .A2(new_n542), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G179), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n545), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n541), .B1(new_n537), .B2(new_n258), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n341), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n539), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(G190), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n572));
  OAI211_X1 g0372(.A(G238), .B(new_n253), .C1(new_n380), .C2(new_n381), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n258), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n266), .A2(G274), .A3(new_n492), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n266), .A2(G250), .A3(new_n501), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n580), .A3(G190), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n258), .B2(new_n575), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n341), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(new_n207), .A3(G33), .A4(G97), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G97), .A2(G107), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n377), .B2(new_n207), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT82), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n252), .A2(new_n590), .A3(new_n207), .A4(G68), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n207), .B(G68), .C1(new_n380), .C2(new_n381), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n279), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n299), .A2(G87), .A3(new_n464), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n320), .A2(new_n303), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n583), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n320), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n299), .A2(new_n464), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT83), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n594), .A2(new_n279), .B1(new_n303), .B2(new_n320), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT83), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n576), .A2(new_n580), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n315), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n582), .A2(new_n346), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n599), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n303), .A2(new_n334), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT25), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n554), .A2(new_n334), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n207), .B(G87), .C1(new_n380), .C2(new_n381), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT22), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT22), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n252), .A2(new_n619), .A3(new_n207), .A4(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n574), .A2(G20), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT23), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n207), .B2(G107), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n334), .A2(KEYINPUT23), .A3(G20), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT24), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT24), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n629), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n616), .B1(new_n631), .B2(new_n279), .ZN(new_n632));
  OAI211_X1 g0432(.A(G257), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n633));
  OAI211_X1 g0433(.A(G250), .B(new_n253), .C1(new_n380), .C2(new_n381), .ZN(new_n634));
  INV_X1    g0434(.A(G33), .ZN(new_n635));
  INV_X1    g0435(.A(G294), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n258), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n503), .A2(G264), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n493), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n315), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n637), .A2(new_n258), .B1(new_n503), .B2(G264), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n346), .A3(new_n493), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT88), .B1(new_n632), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n641), .A2(new_n643), .ZN(new_n646));
  INV_X1    g0446(.A(new_n630), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n629), .B1(new_n621), .B2(new_n626), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n279), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n614), .A2(new_n615), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n640), .A2(G200), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n642), .A2(G190), .A3(new_n493), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n649), .A2(new_n650), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n612), .A2(new_n645), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n463), .A2(new_n529), .A3(new_n571), .A4(new_n657), .ZN(G372));
  OR2_X1    g0458(.A1(new_n398), .A2(new_n349), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n445), .B1(new_n659), .B2(new_n395), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n432), .A2(new_n663), .A3(new_n454), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n432), .B2(new_n454), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n460), .A2(KEYINPUT90), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n448), .A2(new_n663), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n314), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n317), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n605), .A2(new_n595), .A3(new_n597), .A4(new_n601), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n605), .B1(new_n604), .B2(new_n601), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n611), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n599), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n677), .B2(new_n563), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n608), .A2(KEYINPUT89), .A3(new_n315), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT89), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n582), .B2(G169), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n679), .A2(new_n681), .A3(new_n610), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n599), .B1(new_n607), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n567), .A2(new_n568), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n561), .B1(new_n684), .B2(new_n315), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(new_n685), .A3(new_n686), .A4(new_n559), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n607), .A2(new_n682), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n678), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n646), .A2(new_n651), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n516), .B(new_n690), .C1(new_n526), .C2(new_n528), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n673), .A2(new_n674), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n679), .A2(new_n681), .A3(new_n610), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n656), .B(new_n676), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n571), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n672), .B1(new_n463), .B2(new_n698), .ZN(G369));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n513), .A2(new_n515), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n524), .B2(new_n525), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT87), .B1(new_n509), .B2(KEYINPUT21), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n527), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n708));
  INV_X1    g0508(.A(G213), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT93), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n712), .A2(G343), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n704), .B(new_n519), .C1(new_n517), .C2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n516), .B1(new_n526), .B2(new_n528), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n513), .A3(new_n715), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n700), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n645), .A2(new_n653), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n656), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n651), .A2(new_n715), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT94), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n722), .A2(new_n724), .B1(new_n690), .B2(new_n716), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n690), .A2(new_n715), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n722), .A2(new_n724), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n704), .A2(new_n715), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(new_n228), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n586), .A2(new_n587), .A3(new_n471), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n733), .A2(new_n206), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n222), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n733), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT28), .Z(new_n738));
  OAI21_X1  g0538(.A(new_n676), .B1(new_n692), .B2(new_n693), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n739), .B2(new_n563), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n612), .A2(new_n685), .A3(new_n686), .A4(new_n559), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n740), .A2(new_n688), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n645), .A2(new_n653), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n695), .B1(new_n718), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n715), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(KEYINPUT29), .B(new_n715), .C1(new_n689), .C2(new_n696), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n657), .A2(new_n571), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n704), .A3(new_n519), .A4(new_n716), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n642), .A2(new_n582), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n514), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n567), .A3(new_n568), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n753), .A2(new_n567), .A3(KEYINPUT30), .A4(new_n568), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n582), .A2(G179), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n523), .A2(new_n560), .A3(new_n640), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n760), .B2(new_n715), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n700), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n749), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n738), .B1(new_n767), .B2(G1), .ZN(G364));
  NOR2_X1   g0568(.A1(new_n226), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n206), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n733), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n220), .B1(new_n207), .B2(G169), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n276), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n346), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n207), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n780), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n782), .A2(G58), .B1(new_n785), .B2(new_n325), .ZN(new_n786));
  NAND3_X1  g0586(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n276), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n295), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n346), .A2(new_n341), .A3(KEYINPUT98), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT98), .B1(new_n346), .B2(new_n341), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n207), .B1(new_n795), .B2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G97), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n341), .A2(G179), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n779), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G87), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n783), .A2(new_n799), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G107), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n805), .A3(new_n252), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n787), .A2(G190), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G68), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n783), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G159), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n791), .A2(new_n798), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(G294), .ZN(new_n815));
  INV_X1    g0615(.A(G317), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n807), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n819), .B(new_n382), .C1(new_n820), .C2(new_n784), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G326), .B2(new_n788), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n810), .A2(G329), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n800), .B1(new_n781), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G283), .B2(new_n804), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n815), .A2(new_n822), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n778), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT95), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G20), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n777), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n228), .A2(G355), .A3(new_n252), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n246), .A2(new_n261), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n228), .B(new_n382), .C1(G45), .C2(new_n222), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(G116), .B2(new_n228), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n773), .B(new_n829), .C1(new_n833), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n717), .A2(new_n719), .A3(new_n832), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n720), .A2(new_n772), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n717), .A2(new_n700), .A3(new_n719), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  OAI22_X1  g0646(.A1(new_n340), .A2(new_n343), .B1(new_n327), .B2(new_n716), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n349), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n347), .A2(new_n348), .A3(new_n716), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n698), .B2(new_n715), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n344), .A2(new_n349), .A3(new_n716), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n689), .B2(new_n696), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n765), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n772), .B1(new_n855), .B2(new_n765), .ZN(new_n858));
  INV_X1    g0658(.A(new_n831), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n782), .B1(new_n785), .B2(G159), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n788), .A2(G137), .ZN(new_n862));
  INV_X1    g0662(.A(new_n807), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n862), .C1(new_n291), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT34), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n797), .A2(G58), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n252), .B1(new_n803), .B2(new_n352), .C1(new_n295), .C2(new_n800), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G132), .B2(new_n810), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(G283), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n382), .B1(new_n800), .B2(new_n334), .C1(new_n872), .C2(new_n863), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G303), .B2(new_n788), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n810), .A2(G311), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n781), .A2(new_n636), .B1(new_n784), .B2(new_n471), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G87), .B2(new_n804), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n798), .A2(new_n874), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n778), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n778), .A2(new_n831), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT101), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n773), .B(new_n879), .C1(new_n361), .C2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  NOR3_X1   g0684(.A1(new_n222), .A2(new_n210), .A3(new_n421), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n295), .B2(G68), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n886), .A2(new_n206), .A3(G13), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT102), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT36), .ZN(new_n889));
  INV_X1    g0689(.A(new_n549), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n471), .B(new_n221), .C1(new_n890), .C2(KEYINPUT35), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(KEYINPUT35), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  INV_X1    g0694(.A(new_n463), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n751), .A2(new_n763), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT105), .Z(new_n898));
  NAND3_X1  g0698(.A1(new_n425), .A2(new_n430), .A3(new_n283), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n456), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n712), .A2(new_n714), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n460), .A2(new_n449), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n451), .A3(new_n452), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n442), .A2(new_n444), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n432), .A2(new_n901), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n412), .A2(new_n431), .A3(new_n438), .A4(new_n440), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n460), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n900), .A2(new_n454), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n902), .A3(new_n908), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n910), .A2(new_n912), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n906), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n666), .A2(new_n669), .A3(new_n905), .ZN(new_n918));
  INV_X1    g0718(.A(new_n907), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n907), .A2(new_n460), .A3(new_n908), .A4(new_n911), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n909), .B1(new_n667), .B2(new_n668), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n911), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n917), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n371), .A2(new_n715), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n395), .A2(new_n399), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n387), .A2(KEYINPUT14), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n391), .A2(new_n393), .A3(G169), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(new_n346), .C2(new_n391), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n371), .B(new_n715), .C1(new_n930), .C2(new_n398), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n850), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n529), .A2(new_n657), .A3(new_n571), .A4(new_n715), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n760), .A2(new_n715), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT31), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n932), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT40), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n916), .B1(new_n906), .B2(new_n915), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n921), .ZN(new_n943));
  OAI211_X1 g0743(.A(KEYINPUT38), .B(new_n943), .C1(new_n462), .C2(new_n902), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n896), .A3(new_n932), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n700), .B1(new_n898), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n898), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n944), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n927), .A2(new_n931), .ZN(new_n951));
  INV_X1    g0751(.A(new_n849), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n951), .C1(new_n853), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n670), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(new_n901), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(KEYINPUT104), .A3(new_n955), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT39), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n920), .B2(new_n923), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n930), .A2(new_n371), .A3(new_n716), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT39), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n958), .A2(new_n959), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n895), .B1(new_n747), .B2(new_n748), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n672), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n949), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n206), .B2(new_n769), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n949), .A2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n894), .B1(new_n972), .B2(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n228), .A2(new_n382), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n236), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n833), .B1(new_n228), .B2(new_n320), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n772), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n797), .A2(G68), .ZN(new_n979));
  INV_X1    g0779(.A(G159), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n252), .B1(new_n781), .B2(new_n291), .C1(new_n980), .C2(new_n863), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G143), .B2(new_n788), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n810), .A2(G137), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n800), .A2(new_n284), .B1(new_n803), .B2(new_n210), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G50), .B2(new_n785), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n979), .A2(new_n982), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n382), .B1(new_n784), .B2(new_n872), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n781), .A2(new_n824), .B1(new_n803), .B2(new_n468), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G311), .C2(new_n788), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n810), .A2(G317), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n334), .C2(new_n796), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n800), .B2(new_n471), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(new_n863), .C2(new_n636), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT110), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT47), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n777), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n978), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n832), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n715), .A2(new_n598), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n683), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n688), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n743), .A2(new_n570), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n715), .B1(new_n1010), .B2(new_n563), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n728), .A2(new_n729), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n715), .A2(new_n559), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n563), .A2(new_n570), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n685), .A2(new_n559), .A3(new_n715), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT106), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT106), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n728), .A2(new_n729), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1011), .B1(new_n1021), .B2(KEYINPUT42), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT42), .B2(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT107), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1009), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT107), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1008), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n726), .A2(new_n1017), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n733), .B(KEYINPUT41), .Z(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1012), .B1(new_n725), .B2(new_n729), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(new_n720), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n767), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1037), .B(new_n720), .Z(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT108), .B1(new_n1040), .B2(new_n766), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n726), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n730), .A2(new_n1016), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT45), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT44), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n730), .A2(new_n1047), .A3(new_n1016), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n730), .B2(new_n1016), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1042), .B(new_n1043), .C1(new_n1046), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1043), .A2(new_n1042), .ZN(new_n1053));
  AND4_X1   g0853(.A1(new_n1052), .A2(new_n1046), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1039), .B(new_n1041), .C1(new_n1051), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1035), .B1(new_n1055), .B2(new_n767), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1034), .B1(new_n1056), .B2(new_n771), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1033), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1007), .B1(new_n1057), .B2(new_n1058), .ZN(G387));
  OR2_X1    g0859(.A1(new_n725), .A2(new_n1003), .ZN(new_n1060));
  OR3_X1    g0860(.A1(new_n241), .A2(new_n261), .A3(new_n252), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT50), .B1(new_n289), .B2(G50), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n261), .C1(new_n352), .C2(new_n361), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n382), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n734), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n732), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n833), .B1(new_n334), .B2(new_n228), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n772), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n797), .A2(new_n600), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n252), .B1(new_n803), .B2(new_n468), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n789), .A2(new_n980), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n288), .C2(new_n807), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n810), .A2(G150), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n295), .A2(new_n781), .B1(new_n800), .B2(new_n210), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G68), .B2(new_n785), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n810), .A2(G326), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n252), .B1(new_n804), .B2(G116), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G317), .A2(new_n782), .B1(new_n785), .B2(G303), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n789), .B2(new_n825), .C1(new_n820), .C2(new_n863), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT48), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n796), .A2(new_n872), .B1(new_n636), .B2(new_n800), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(KEYINPUT111), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(KEYINPUT111), .B2(new_n1084), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT49), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1079), .B(new_n1080), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1078), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1070), .B1(new_n1090), .B2(new_n777), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1038), .A2(new_n771), .B1(new_n1060), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n733), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1094), .A2(new_n1095), .B1(new_n767), .B2(new_n1038), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(G393));
  NOR2_X1   g0898(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n733), .A3(new_n1055), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n771), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n833), .B1(new_n468), .B2(new_n228), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n250), .A2(new_n975), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n772), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n800), .A2(new_n872), .B1(new_n784), .B2(new_n636), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n805), .A2(new_n382), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G303), .C2(new_n807), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n789), .A2(new_n816), .B1(new_n781), .B2(new_n820), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT52), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n797), .A2(G116), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n810), .A2(G322), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n782), .A2(G159), .B1(G150), .B2(new_n788), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT113), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT51), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n289), .A2(new_n784), .B1(new_n800), .B2(new_n352), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n382), .B(new_n1118), .C1(G87), .C2(new_n804), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n797), .A2(G77), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n810), .A2(G143), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n807), .A2(G50), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1114), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1106), .B1(new_n1124), .B2(new_n777), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1016), .B2(new_n1003), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1102), .A2(new_n1103), .A3(new_n1126), .ZN(G390));
  AOI21_X1  g0927(.A(new_n773), .B1(new_n881), .B2(new_n289), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT117), .Z(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n789), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n801), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G137), .C2(new_n807), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n797), .A2(G159), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n810), .A2(G125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n784), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n252), .B1(new_n803), .B2(new_n295), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(G132), .C2(new_n782), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n802), .B(new_n382), .C1(new_n872), .C2(new_n789), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G107), .B2(new_n807), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n810), .A2(G294), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n781), .A2(new_n471), .B1(new_n803), .B2(new_n352), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G97), .B2(new_n785), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1120), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n962), .A2(new_n965), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1129), .B1(new_n778), .B2(new_n1148), .C1(new_n1150), .C2(new_n831), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n850), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n1153), .C1(new_n933), .C2(new_n938), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n951), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n951), .B1(new_n853), .B2(new_n952), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n962), .A2(new_n965), .B1(new_n1157), .B2(new_n963), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n963), .B1(new_n961), .B2(new_n917), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n683), .A2(new_n563), .A3(new_n570), .A4(new_n656), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n704), .B2(new_n721), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n740), .A2(new_n688), .A3(new_n741), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n716), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n848), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n849), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1159), .B1(new_n1165), .B2(new_n951), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1156), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n852), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n952), .B1(new_n697), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n963), .B1(new_n1169), .B2(new_n1155), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1149), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n924), .A2(new_n916), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n964), .B1(new_n1172), .B2(new_n944), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n952), .B1(new_n745), .B2(new_n848), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n1155), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n764), .A2(new_n1153), .A3(new_n951), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1167), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n770), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1152), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1169), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n951), .B1(new_n764), .B2(new_n1153), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1156), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n895), .A2(new_n764), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n968), .A2(new_n672), .A3(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1167), .A2(new_n1186), .A3(new_n1177), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n733), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT114), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT114), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1192), .A3(new_n733), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1178), .A2(KEYINPUT115), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT115), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1167), .A2(new_n1196), .A3(new_n1177), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT116), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1189), .A2(new_n1192), .A3(new_n733), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1192), .B1(new_n1189), .B2(new_n733), .ZN(new_n1202));
  OAI211_X1 g1002(.A(KEYINPUT116), .B(new_n1199), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1180), .B1(new_n1200), .B2(new_n1204), .ZN(G378));
  OAI21_X1  g1005(.A(new_n772), .B1(new_n880), .B2(G50), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT119), .Z(new_n1207));
  NOR2_X1   g1007(.A1(new_n252), .A2(G41), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G50), .B(new_n1208), .C1(new_n635), .C2(new_n260), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n600), .A2(new_n785), .B1(new_n804), .B2(G58), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n334), .B2(new_n781), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G283), .B2(new_n810), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1208), .B1(new_n800), .B2(new_n210), .C1(new_n468), .C2(new_n863), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n788), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n979), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1130), .A2(new_n781), .B1(new_n800), .B2(new_n1137), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G137), .B2(new_n785), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n807), .A2(G132), .B1(new_n788), .B2(G125), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n291), .C2(new_n796), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n635), .B(new_n260), .C1(new_n803), .C2(new_n980), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n810), .B2(G124), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1222), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1207), .B1(new_n1227), .B2(new_n777), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n901), .A2(new_n305), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n318), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n314), .A2(new_n317), .A3(new_n1229), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1228), .B1(new_n1237), .B2(new_n831), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n947), .B2(G330), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n700), .B(new_n1236), .C1(new_n940), .C2(new_n946), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n967), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n896), .B(new_n932), .C1(new_n961), .C2(new_n917), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n939), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(KEYINPUT40), .A2(new_n1243), .B1(new_n1244), .B2(new_n945), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1236), .B1(new_n1245), .B2(new_n700), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1150), .A2(new_n964), .B1(new_n956), .B2(new_n957), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n947), .A2(G330), .A3(new_n1237), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n959), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1239), .B1(new_n1250), .B2(new_n771), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1249), .A2(new_n1242), .B1(new_n1189), .B2(new_n1188), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n733), .B1(new_n1252), .B2(KEYINPUT57), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1189), .A2(new_n1188), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1250), .A2(KEYINPUT57), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1251), .B1(new_n1253), .B2(new_n1255), .ZN(G375));
  INV_X1    g1056(.A(new_n1035), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n968), .A2(new_n672), .A3(new_n1187), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1198), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1155), .A2(new_n859), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G137), .A2(new_n782), .B1(new_n785), .B2(G150), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n980), .B2(new_n800), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G128), .B2(new_n810), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n252), .B1(new_n803), .B2(new_n284), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n863), .A2(new_n1137), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(G132), .C2(new_n788), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1264), .B(new_n1267), .C1(new_n295), .C2(new_n796), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n800), .A2(new_n468), .B1(new_n784), .B2(new_n334), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n863), .A2(new_n471), .B1(new_n789), .B2(new_n636), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G283), .C2(new_n782), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n810), .A2(G303), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n382), .B1(new_n803), .B2(new_n361), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT121), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1071), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n778), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n773), .B(new_n1276), .C1(new_n352), .C2(new_n881), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1186), .A2(new_n771), .B1(new_n1261), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1260), .A2(new_n1278), .ZN(G381));
  INV_X1    g1079(.A(G390), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n883), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(new_n1281), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1282));
  INV_X1    g1082(.A(G387), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1199), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n1180), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1286), .ZN(G407));
  NOR2_X1   g1087(.A1(new_n709), .A2(G343), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G407), .A2(G213), .A3(new_n1289), .ZN(G409));
  NAND2_X1  g1090(.A1(new_n1288), .A2(G2897), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1258), .A2(new_n1183), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n733), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1198), .A2(KEYINPUT60), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1259), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1278), .ZN(new_n1297));
  OR3_X1    g1097(.A1(new_n1296), .A2(new_n883), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n883), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT122), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1292), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1302), .A2(new_n1292), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT123), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G378), .A2(new_n1284), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1250), .A2(new_n771), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1238), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1286), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1288), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT123), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1303), .A2(new_n1304), .A3(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1306), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G387), .A2(new_n1280), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(G393), .B(new_n845), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1033), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1321), .B(new_n1034), .C1(new_n771), .C2(new_n1056), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1007), .A3(G390), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1317), .A2(new_n1318), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1318), .B1(new_n1317), .B2(new_n1323), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT61), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1288), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT116), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1285), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1203), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G375), .B1(new_n1332), .B2(new_n1180), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1286), .A2(new_n1310), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1327), .B(new_n1329), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1329), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1316), .A2(new_n1326), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT124), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1335), .A2(new_n1340), .A3(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1312), .B2(new_n1305), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT62), .B1(new_n1335), .B2(new_n1340), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1339), .B1(new_n1345), .B2(new_n1346), .ZN(G405));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1348), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1318), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(G387), .A2(new_n1280), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G390), .B1(new_n1322), .B2(new_n1007), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1350), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1317), .A2(new_n1323), .A3(new_n1318), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1353), .A2(KEYINPUT127), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1349), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G375), .A2(new_n1286), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1329), .A2(KEYINPUT126), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT126), .B1(new_n1329), .B2(KEYINPUT125), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n1307), .B(new_n1357), .C1(new_n1358), .C2(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1333), .B1(G375), .B2(new_n1286), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1360), .B1(new_n1361), .B2(new_n1359), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1356), .B(new_n1362), .ZN(G402));
endmodule


