

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n724), .ZN(n698) );
  NAND2_X1 U549 ( .A1(n761), .A2(n759), .ZN(n724) );
  NOR2_X1 U550 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U551 ( .A1(n868), .A2(G137), .ZN(n527) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n521), .ZN(n531) );
  AND2_X1 U553 ( .A1(n791), .A2(n804), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n758), .A2(n757), .ZN(n515) );
  AND2_X1 U555 ( .A1(n698), .A2(G1996), .ZN(n680) );
  INV_X1 U556 ( .A(KEYINPUT91), .ZN(n710) );
  XNOR2_X1 U557 ( .A(n710), .B(KEYINPUT31), .ZN(n711) );
  XNOR2_X1 U558 ( .A(n712), .B(n711), .ZN(n713) );
  INV_X1 U559 ( .A(KEYINPUT93), .ZN(n719) );
  NAND2_X1 U560 ( .A1(G8), .A2(n724), .ZN(n752) );
  XNOR2_X1 U561 ( .A(n674), .B(KEYINPUT83), .ZN(n759) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U563 ( .A1(G651), .A2(n643), .ZN(n638) );
  NOR2_X1 U564 ( .A1(n525), .A2(n524), .ZN(G164) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XNOR2_X2 U566 ( .A(n517), .B(n516), .ZN(n868) );
  NAND2_X1 U567 ( .A1(G138), .A2(n868), .ZN(n518) );
  XNOR2_X1 U568 ( .A(n518), .B(KEYINPUT82), .ZN(n520) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n862) );
  NAND2_X1 U570 ( .A1(n862), .A2(G114), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n525) );
  XNOR2_X1 U572 ( .A(G2104), .B(KEYINPUT65), .ZN(n521) );
  NAND2_X1 U573 ( .A1(G102), .A2(n531), .ZN(n523) );
  AND2_X1 U574 ( .A1(n521), .A2(G2105), .ZN(n864) );
  NAND2_X1 U575 ( .A1(G126), .A2(n864), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G113), .A2(n862), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(n528), .ZN(n530) );
  AND2_X1 U580 ( .A1(n864), .A2(G125), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n673) );
  NAND2_X1 U582 ( .A1(G101), .A2(n531), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n532), .Z(n671) );
  AND2_X1 U584 ( .A1(n673), .A2(n671), .ZN(G160) );
  AND2_X1 U585 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U586 ( .A(G132), .ZN(G219) );
  INV_X1 U587 ( .A(G82), .ZN(G220) );
  INV_X1 U588 ( .A(G57), .ZN(G237) );
  INV_X1 U589 ( .A(G120), .ZN(G236) );
  INV_X1 U590 ( .A(G651), .ZN(n536) );
  NOR2_X1 U591 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n533), .Z(n642) );
  NAND2_X1 U593 ( .A1(G64), .A2(n642), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  NAND2_X1 U595 ( .A1(G52), .A2(n638), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n543) );
  OR2_X1 U597 ( .A1(n536), .A2(n643), .ZN(n537) );
  XNOR2_X1 U598 ( .A(KEYINPUT67), .B(n537), .ZN(n631) );
  NAND2_X1 U599 ( .A1(n631), .A2(G77), .ZN(n540) );
  NOR2_X1 U600 ( .A1(G543), .A2(G651), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT64), .ZN(n628) );
  NAND2_X1 U602 ( .A1(G90), .A2(n628), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(G171) );
  NAND2_X1 U606 ( .A1(G7), .A2(G661), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U608 ( .A(G223), .ZN(n810) );
  NAND2_X1 U609 ( .A1(n810), .A2(G567), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT11), .B(n545), .Z(G234) );
  NAND2_X1 U611 ( .A1(G81), .A2(n628), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT12), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G68), .A2(n631), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT13), .B(n549), .Z(n553) );
  NAND2_X1 U616 ( .A1(G56), .A2(n642), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT69), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT14), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n638), .A2(G43), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n942) );
  INV_X1 U622 ( .A(G860), .ZN(n606) );
  OR2_X1 U623 ( .A1(n942), .A2(n606), .ZN(G153) );
  INV_X1 U624 ( .A(G171), .ZN(G301) );
  NAND2_X1 U625 ( .A1(G301), .A2(G868), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n556), .B(KEYINPUT70), .ZN(n565) );
  INV_X1 U627 ( .A(G868), .ZN(n654) );
  NAND2_X1 U628 ( .A1(G66), .A2(n642), .ZN(n558) );
  NAND2_X1 U629 ( .A1(G54), .A2(n638), .ZN(n557) );
  NAND2_X1 U630 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n631), .A2(G79), .ZN(n560) );
  NAND2_X1 U632 ( .A1(G92), .A2(n628), .ZN(n559) );
  NAND2_X1 U633 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n563), .B(KEYINPUT15), .ZN(n925) );
  NAND2_X1 U636 ( .A1(n654), .A2(n925), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(G284) );
  XNOR2_X1 U638 ( .A(KEYINPUT6), .B(KEYINPUT72), .ZN(n569) );
  NAND2_X1 U639 ( .A1(G63), .A2(n642), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G51), .A2(n638), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U642 ( .A(n569), .B(n568), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n628), .A2(G89), .ZN(n570) );
  XOR2_X1 U644 ( .A(KEYINPUT71), .B(n570), .Z(n571) );
  XNOR2_X1 U645 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U646 ( .A1(G76), .A2(n631), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U648 ( .A(KEYINPUT5), .B(n574), .Z(n575) );
  NOR2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U650 ( .A(KEYINPUT73), .B(KEYINPUT7), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n578), .B(n577), .ZN(G168) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(n579) );
  XNOR2_X1 U653 ( .A(KEYINPUT74), .B(n579), .ZN(G286) );
  NAND2_X1 U654 ( .A1(G65), .A2(n642), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G53), .A2(n638), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n631), .A2(G78), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G91), .A2(n628), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n934) );
  XOR2_X1 U661 ( .A(n934), .B(KEYINPUT68), .Z(G299) );
  NAND2_X1 U662 ( .A1(G868), .A2(G286), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G299), .A2(n654), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n606), .A2(G559), .ZN(n588) );
  INV_X1 U666 ( .A(n925), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n588), .A2(n604), .ZN(n589) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n942), .ZN(n592) );
  NAND2_X1 U670 ( .A1(G868), .A2(n604), .ZN(n590) );
  NOR2_X1 U671 ( .A1(G559), .A2(n590), .ZN(n591) );
  NOR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G111), .A2(n862), .ZN(n594) );
  NAND2_X1 U674 ( .A1(G99), .A2(n531), .ZN(n593) );
  NAND2_X1 U675 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U676 ( .A(KEYINPUT76), .B(n595), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n864), .A2(G123), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U679 ( .A1(G135), .A2(n868), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U681 ( .A(KEYINPUT75), .B(n599), .Z(n600) );
  NOR2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n963) );
  XNOR2_X1 U683 ( .A(G2096), .B(n963), .ZN(n603) );
  INV_X1 U684 ( .A(G2100), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G559), .A2(n604), .ZN(n605) );
  XOR2_X1 U687 ( .A(n942), .B(n605), .Z(n652) );
  NAND2_X1 U688 ( .A1(n606), .A2(n652), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G80), .A2(n631), .ZN(n608) );
  NAND2_X1 U690 ( .A1(G67), .A2(n642), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U692 ( .A1(G93), .A2(n628), .ZN(n609) );
  XNOR2_X1 U693 ( .A(KEYINPUT77), .B(n609), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n638), .A2(G55), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n655) );
  XNOR2_X1 U697 ( .A(n614), .B(n655), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G75), .A2(n631), .ZN(n616) );
  NAND2_X1 U699 ( .A1(G62), .A2(n642), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G88), .A2(n628), .ZN(n617) );
  XNOR2_X1 U702 ( .A(KEYINPUT79), .B(n617), .ZN(n618) );
  NOR2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n638), .A2(G50), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(G303) );
  INV_X1 U706 ( .A(G303), .ZN(G166) );
  AND2_X1 U707 ( .A1(n631), .A2(G72), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n638), .A2(G47), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G85), .A2(n628), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n642), .A2(G60), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G48), .A2(n638), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n642), .A2(G61), .ZN(n630) );
  NAND2_X1 U716 ( .A1(G86), .A2(n628), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n631), .A2(G73), .ZN(n632) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U722 ( .A(n637), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G49), .A2(n638), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n643), .A2(G87), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G288) );
  XNOR2_X1 U729 ( .A(G166), .B(G299), .ZN(n647) );
  XNOR2_X1 U730 ( .A(G290), .B(G305), .ZN(n646) );
  XNOR2_X1 U731 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U732 ( .A(n648), .B(G288), .ZN(n651) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n649) );
  XNOR2_X1 U734 ( .A(n649), .B(n655), .ZN(n650) );
  XNOR2_X1 U735 ( .A(n651), .B(n650), .ZN(n880) );
  XOR2_X1 U736 ( .A(n880), .B(n652), .Z(n653) );
  NOR2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n657) );
  NOR2_X1 U738 ( .A1(G868), .A2(n655), .ZN(n656) );
  NOR2_X1 U739 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G236), .A2(G237), .ZN(n662) );
  NAND2_X1 U747 ( .A1(G69), .A2(n662), .ZN(n663) );
  XNOR2_X1 U748 ( .A(KEYINPUT81), .B(n663), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n664), .A2(G108), .ZN(n814) );
  NAND2_X1 U750 ( .A1(n814), .A2(G567), .ZN(n669) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n665), .Z(n666) );
  NOR2_X1 U753 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U754 ( .A1(G96), .A2(n667), .ZN(n815) );
  NAND2_X1 U755 ( .A1(n815), .A2(G2106), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n816) );
  NAND2_X1 U757 ( .A1(G661), .A2(G483), .ZN(n670) );
  NOR2_X1 U758 ( .A1(n816), .A2(n670), .ZN(n813) );
  NAND2_X1 U759 ( .A1(n813), .A2(G36), .ZN(G176) );
  XNOR2_X1 U760 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n809) );
  NOR2_X1 U761 ( .A1(G164), .A2(G1384), .ZN(n761) );
  AND2_X1 U762 ( .A1(G40), .A2(n671), .ZN(n672) );
  NAND2_X1 U763 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n931) );
  NAND2_X1 U765 ( .A1(n931), .A2(KEYINPUT33), .ZN(n675) );
  NOR2_X1 U766 ( .A1(n752), .A2(n675), .ZN(n742) );
  NOR2_X1 U767 ( .A1(G2084), .A2(n724), .ZN(n703) );
  NAND2_X1 U768 ( .A1(G8), .A2(n703), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n698), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U770 ( .A(n676), .B(KEYINPUT27), .ZN(n678) );
  AND2_X1 U771 ( .A1(G1956), .A2(n724), .ZN(n677) );
  NOR2_X1 U772 ( .A1(n678), .A2(n677), .ZN(n691) );
  NOR2_X1 U773 ( .A1(n934), .A2(n691), .ZN(n679) );
  XOR2_X1 U774 ( .A(n679), .B(KEYINPUT28), .Z(n695) );
  XOR2_X1 U775 ( .A(n680), .B(KEYINPUT26), .Z(n682) );
  NAND2_X1 U776 ( .A1(n724), .A2(G1341), .ZN(n681) );
  NAND2_X1 U777 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U778 ( .A1(n942), .A2(n683), .ZN(n687) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n724), .ZN(n685) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n698), .ZN(n684) );
  NAND2_X1 U781 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U782 ( .A1(n925), .A2(n688), .ZN(n686) );
  OR2_X1 U783 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n925), .A2(n688), .ZN(n689) );
  NAND2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n934), .A2(n691), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT29), .ZN(n702) );
  XOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .Z(n901) );
  NOR2_X1 U791 ( .A1(n901), .A2(n724), .ZN(n697) );
  XNOR2_X1 U792 ( .A(n697), .B(KEYINPUT90), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n698), .A2(G1961), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n707) );
  NOR2_X1 U795 ( .A1(G301), .A2(n707), .ZN(n701) );
  NOR2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n714) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n752), .ZN(n717) );
  NOR2_X1 U798 ( .A1(n703), .A2(n717), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n704), .A2(G8), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT30), .ZN(n706) );
  NOR2_X1 U801 ( .A1(G168), .A2(n706), .ZN(n709) );
  AND2_X1 U802 ( .A1(G301), .A2(n707), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n716) );
  INV_X1 U805 ( .A(KEYINPUT92), .ZN(n715) );
  XNOR2_X1 U806 ( .A(n716), .B(n715), .ZN(n723) );
  INV_X1 U807 ( .A(n723), .ZN(n718) );
  XNOR2_X1 U808 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n733) );
  NAND2_X1 U810 ( .A1(n723), .A2(G286), .ZN(n729) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n752), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n727), .A2(G303), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U816 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U817 ( .A(n731), .B(KEYINPUT32), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n749) );
  NOR2_X1 U819 ( .A1(G1971), .A2(G303), .ZN(n734) );
  XNOR2_X1 U820 ( .A(KEYINPUT94), .B(n734), .ZN(n735) );
  NOR2_X1 U821 ( .A1(n931), .A2(n735), .ZN(n736) );
  XOR2_X1 U822 ( .A(KEYINPUT95), .B(n736), .Z(n737) );
  NAND2_X1 U823 ( .A1(n749), .A2(n737), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U825 ( .A1(n738), .A2(n932), .ZN(n739) );
  NOR2_X1 U826 ( .A1(n752), .A2(n739), .ZN(n740) );
  NOR2_X1 U827 ( .A1(KEYINPUT33), .A2(n740), .ZN(n741) );
  NOR2_X1 U828 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U829 ( .A(G1981), .B(G305), .Z(n928) );
  NAND2_X1 U830 ( .A1(n743), .A2(n928), .ZN(n758) );
  NOR2_X1 U831 ( .A1(G1981), .A2(G305), .ZN(n744) );
  XNOR2_X1 U832 ( .A(KEYINPUT24), .B(n744), .ZN(n745) );
  XNOR2_X1 U833 ( .A(KEYINPUT89), .B(n745), .ZN(n746) );
  OR2_X1 U834 ( .A1(n752), .A2(n746), .ZN(n756) );
  INV_X1 U835 ( .A(KEYINPUT97), .ZN(n754) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n747) );
  XNOR2_X1 U837 ( .A(n747), .B(KEYINPUT96), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n748), .A2(G8), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n754), .B(n753), .ZN(n755) );
  AND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n757) );
  INV_X1 U843 ( .A(n759), .ZN(n760) );
  NOR2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n804) );
  NAND2_X1 U845 ( .A1(G140), .A2(n868), .ZN(n763) );
  NAND2_X1 U846 ( .A1(G104), .A2(n531), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U848 ( .A(KEYINPUT34), .B(n764), .ZN(n769) );
  NAND2_X1 U849 ( .A1(G116), .A2(n862), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G128), .A2(n864), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U852 ( .A(KEYINPUT35), .B(n767), .Z(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n770), .ZN(n853) );
  XNOR2_X1 U855 ( .A(KEYINPUT37), .B(G2067), .ZN(n802) );
  NOR2_X1 U856 ( .A1(n853), .A2(n802), .ZN(n964) );
  NAND2_X1 U857 ( .A1(n804), .A2(n964), .ZN(n771) );
  XOR2_X1 U858 ( .A(KEYINPUT84), .B(n771), .Z(n800) );
  NAND2_X1 U859 ( .A1(G131), .A2(n868), .ZN(n772) );
  XNOR2_X1 U860 ( .A(n772), .B(KEYINPUT86), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G95), .A2(n531), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G119), .A2(n864), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G107), .A2(n862), .ZN(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT85), .B(n775), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n854) );
  NAND2_X1 U868 ( .A1(G1991), .A2(n854), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT87), .ZN(n790) );
  NAND2_X1 U870 ( .A1(G117), .A2(n862), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G129), .A2(n864), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n531), .A2(G105), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(KEYINPUT88), .B(n786), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G141), .A2(n868), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n875) );
  AND2_X1 U879 ( .A1(G1996), .A2(n875), .ZN(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n955) );
  XOR2_X1 U881 ( .A(G1986), .B(G290), .Z(n924) );
  NAND2_X1 U882 ( .A1(n955), .A2(n924), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n800), .A2(n514), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n515), .A2(n792), .ZN(n807) );
  NOR2_X1 U885 ( .A1(G1991), .A2(n854), .ZN(n962) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n793) );
  NOR2_X1 U887 ( .A1(n962), .A2(n793), .ZN(n795) );
  INV_X1 U888 ( .A(n955), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n797) );
  NOR2_X1 U890 ( .A1(n875), .A2(G1996), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n796), .B(KEYINPUT98), .ZN(n952) );
  NOR2_X1 U892 ( .A1(n797), .A2(n952), .ZN(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT39), .B(n798), .Z(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT99), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n853), .A2(n802), .ZN(n954) );
  NAND2_X1 U897 ( .A1(n803), .A2(n954), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U900 ( .A(n809), .B(n808), .ZN(G329) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n810), .ZN(G217) );
  AND2_X1 U902 ( .A1(G15), .A2(G2), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G661), .A2(n811), .ZN(G259) );
  NAND2_X1 U904 ( .A1(G3), .A2(G1), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(G188) );
  XOR2_X1 U906 ( .A(G108), .B(KEYINPUT110), .Z(G238) );
  INV_X1 U908 ( .A(G96), .ZN(G221) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(G325) );
  INV_X1 U910 ( .A(G325), .ZN(G261) );
  INV_X1 U911 ( .A(n816), .ZN(G319) );
  XOR2_X1 U912 ( .A(G2096), .B(KEYINPUT43), .Z(n818) );
  XNOR2_X1 U913 ( .A(G2090), .B(KEYINPUT102), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U915 ( .A(n819), .B(G2678), .Z(n821) );
  XNOR2_X1 U916 ( .A(G2067), .B(G2072), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n821), .B(n820), .ZN(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT42), .B(G2100), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2084), .B(G2078), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n825), .B(n824), .ZN(G227) );
  XOR2_X1 U922 ( .A(G1956), .B(G1966), .Z(n827) );
  XNOR2_X1 U923 ( .A(G1986), .B(G1981), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U925 ( .A(G1971), .B(G1976), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U929 ( .A(KEYINPUT103), .B(G2474), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n835) );
  XOR2_X1 U931 ( .A(G1961), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(G229) );
  NAND2_X1 U933 ( .A1(G124), .A2(n864), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT44), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n862), .A2(G112), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G136), .A2(n868), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G100), .A2(n531), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(G162) );
  NAND2_X1 U941 ( .A1(G142), .A2(n868), .ZN(n844) );
  NAND2_X1 U942 ( .A1(G106), .A2(n531), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n845), .B(KEYINPUT45), .ZN(n847) );
  NAND2_X1 U945 ( .A1(G130), .A2(n864), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n862), .A2(G118), .ZN(n848) );
  XOR2_X1 U948 ( .A(KEYINPUT104), .B(n848), .Z(n849) );
  NOR2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(G160), .B(n851), .Z(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n858) );
  XNOR2_X1 U952 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n854), .B(KEYINPUT108), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U956 ( .A(G164), .B(G162), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(n861), .B(n963), .Z(n877) );
  NAND2_X1 U959 ( .A1(n862), .A2(G115), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n863), .B(KEYINPUT106), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G127), .A2(n864), .ZN(n865) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U963 ( .A(n867), .B(KEYINPUT47), .ZN(n870) );
  NAND2_X1 U964 ( .A1(G139), .A2(n868), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G103), .A2(n531), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT105), .B(n871), .ZN(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n874), .Z(n956) );
  XOR2_X1 U970 ( .A(n875), .B(n956), .Z(n876) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U972 ( .A1(G37), .A2(n878), .ZN(n879) );
  XOR2_X1 U973 ( .A(KEYINPUT109), .B(n879), .Z(G395) );
  XNOR2_X1 U974 ( .A(n880), .B(n942), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n881), .B(G286), .ZN(n883) );
  XNOR2_X1 U976 ( .A(n925), .B(G171), .ZN(n882) );
  XNOR2_X1 U977 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U978 ( .A1(G37), .A2(n884), .ZN(G397) );
  XOR2_X1 U979 ( .A(G2454), .B(G2430), .Z(n886) );
  XNOR2_X1 U980 ( .A(G2451), .B(G2446), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n893) );
  XOR2_X1 U982 ( .A(G2443), .B(G2427), .Z(n888) );
  XNOR2_X1 U983 ( .A(G2438), .B(KEYINPUT101), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(G2435), .Z(n891) );
  XNOR2_X1 U986 ( .A(G1341), .B(G1348), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n894), .A2(G14), .ZN(n900) );
  NAND2_X1 U990 ( .A1(G319), .A2(n900), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT49), .B(n895), .ZN(n896) );
  NOR2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G395), .A2(G397), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(G225) );
  INV_X1 U996 ( .A(G225), .ZN(G308) );
  INV_X1 U997 ( .A(G69), .ZN(G235) );
  INV_X1 U998 ( .A(n900), .ZN(G401) );
  XNOR2_X1 U999 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1011) );
  XOR2_X1 U1000 ( .A(G2090), .B(G35), .Z(n915) );
  XNOR2_X1 U1001 ( .A(G1996), .B(G32), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G27), .B(n901), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n911) );
  XOR2_X1 U1004 ( .A(G1991), .B(G25), .Z(n904) );
  NAND2_X1 U1005 ( .A1(n904), .A2(G28), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G26), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(G2072), .B(G33), .ZN(n905) );
  NOR2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n907), .B(KEYINPUT113), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(KEYINPUT114), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(KEYINPUT53), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(G34), .B(G2084), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT54), .B(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT115), .B(n919), .Z(n920) );
  NOR2_X1 U1019 ( .A1(G29), .A2(n920), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT55), .B(n921), .Z(n1009) );
  XNOR2_X1 U1021 ( .A(G1961), .B(KEYINPUT117), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(G301), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(G1348), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n946) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G168), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT57), .ZN(n941) );
  INV_X1 U1029 ( .A(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(G166), .B(G1971), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n934), .B(G1956), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT118), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G1341), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n947), .B(KEYINPUT116), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(KEYINPUT119), .ZN(n1006) );
  XOR2_X1 U1044 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT51), .B(n953), .Z(n973) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n971) );
  XOR2_X1 U1048 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(KEYINPUT112), .B(n959), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n960), .B(KEYINPUT50), .ZN(n969) );
  XOR2_X1 U1053 ( .A(G160), .B(G2084), .Z(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n966) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(KEYINPUT111), .B(n967), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1060 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1061 ( .A(n974), .B(KEYINPUT52), .ZN(n975) );
  NAND2_X1 U1062 ( .A1(n975), .A2(G29), .ZN(n1004) );
  XOR2_X1 U1063 ( .A(G16), .B(KEYINPUT120), .Z(n1002) );
  XOR2_X1 U1064 ( .A(G1986), .B(G24), .Z(n978) );
  XOR2_X1 U1065 ( .A(G22), .B(KEYINPUT124), .Z(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(G1971), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1068 ( .A(KEYINPUT125), .B(G1976), .Z(n979) );
  XNOR2_X1 U1069 ( .A(G23), .B(n979), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1071 ( .A(KEYINPUT58), .B(n982), .Z(n999) );
  XOR2_X1 U1072 ( .A(G1961), .B(G5), .Z(n994) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G19), .B(G1341), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT121), .B(n985), .Z(n989) );
  XNOR2_X1 U1077 ( .A(KEYINPUT59), .B(G4), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT122), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n987), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G20), .B(G1956), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n992), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G21), .B(G1966), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT123), .B(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(KEYINPUT61), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(G11), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1012), .ZN(G150) );
  INV_X1 U1097 ( .A(G150), .ZN(G311) );
endmodule

