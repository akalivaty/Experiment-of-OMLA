

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(KEYINPUT1), .B(n545), .ZN(n802) );
  AND2_X2 U555 ( .A1(n527), .A2(G2104), .ZN(n892) );
  NOR2_X1 U556 ( .A1(n664), .A2(n786), .ZN(n658) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n633) );
  OR2_X1 U558 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U559 ( .A1(n737), .A2(n736), .ZN(n739) );
  NOR2_X1 U560 ( .A1(n990), .A2(n648), .ZN(n649) );
  XNOR2_X1 U561 ( .A(n675), .B(KEYINPUT91), .ZN(n659) );
  INV_X1 U562 ( .A(n659), .ZN(n677) );
  INV_X1 U563 ( .A(KEYINPUT103), .ZN(n738) );
  XNOR2_X1 U564 ( .A(n739), .B(n738), .ZN(n740) );
  INV_X1 U565 ( .A(G651), .ZN(n543) );
  NAND2_X1 U566 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U567 ( .A1(G543), .A2(G651), .ZN(n805) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n527), .ZN(n889) );
  AND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U570 ( .A1(n888), .A2(G114), .ZN(n522) );
  XNOR2_X1 U571 ( .A(n522), .B(KEYINPUT84), .ZN(n526) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U574 ( .A(n524), .B(n523), .ZN(n591) );
  NAND2_X1 U575 ( .A1(G138), .A2(n591), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n531) );
  INV_X1 U577 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G102), .A2(n892), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G126), .A2(n889), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U582 ( .A1(n888), .A2(G113), .ZN(n534) );
  NAND2_X1 U583 ( .A1(G101), .A2(n892), .ZN(n532) );
  XOR2_X1 U584 ( .A(n532), .B(KEYINPUT23), .Z(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G137), .A2(n591), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G125), .A2(n889), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U589 ( .A1(n538), .A2(n537), .ZN(G160) );
  NAND2_X1 U590 ( .A1(G90), .A2(n805), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n567) );
  NOR2_X1 U592 ( .A1(n567), .A2(n543), .ZN(n806) );
  NAND2_X1 U593 ( .A1(G77), .A2(n806), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT9), .B(n541), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n567), .A2(G651), .ZN(n542) );
  XNOR2_X1 U597 ( .A(KEYINPUT64), .B(n542), .ZN(n801) );
  NAND2_X1 U598 ( .A1(n801), .A2(G52), .ZN(n547) );
  NOR2_X1 U599 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U600 ( .A(KEYINPUT66), .B(n544), .Z(n545) );
  NAND2_X1 U601 ( .A1(n802), .A2(G64), .ZN(n546) );
  AND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(G301) );
  INV_X1 U604 ( .A(G301), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n805), .A2(G89), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G76), .A2(n806), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G51), .A2(n801), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT72), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G63), .A2(n802), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U617 ( .A1(G88), .A2(n805), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G75), .A2(n806), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G50), .A2(n801), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G62), .A2(n802), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U623 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U626 ( .A1(G87), .A2(n567), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G651), .A2(G74), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G49), .A2(n801), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U630 ( .A1(n802), .A2(n570), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n573), .B(KEYINPUT78), .ZN(G288) );
  NAND2_X1 U633 ( .A1(n805), .A2(G86), .ZN(n580) );
  NAND2_X1 U634 ( .A1(G48), .A2(n801), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G61), .A2(n802), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n806), .A2(G73), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U641 ( .A(KEYINPUT79), .B(n581), .Z(G305) );
  NAND2_X1 U642 ( .A1(G85), .A2(n805), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G72), .A2(n806), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G47), .A2(n801), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G60), .A2(n802), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT67), .B(n586), .Z(n587) );
  NOR2_X1 U649 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U650 ( .A(KEYINPUT68), .B(n589), .Z(G290) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n620) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n619) );
  NOR2_X1 U653 ( .A1(n620), .A2(n619), .ZN(n757) );
  NAND2_X1 U654 ( .A1(n892), .A2(G104), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(KEYINPUT86), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G140), .A2(n591), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(KEYINPUT34), .B(n594), .ZN(n599) );
  NAND2_X1 U659 ( .A1(G116), .A2(n888), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G128), .A2(n889), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U662 ( .A(KEYINPUT35), .B(n597), .Z(n598) );
  NOR2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(KEYINPUT36), .B(n600), .ZN(n903) );
  XNOR2_X1 U665 ( .A(G2067), .B(KEYINPUT37), .ZN(n755) );
  NOR2_X1 U666 ( .A1(n903), .A2(n755), .ZN(n930) );
  NAND2_X1 U667 ( .A1(n757), .A2(n930), .ZN(n752) );
  NAND2_X1 U668 ( .A1(n889), .A2(G119), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G131), .A2(n591), .ZN(n601) );
  XOR2_X1 U670 ( .A(KEYINPUT87), .B(n601), .Z(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G107), .A2(n888), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G95), .A2(n892), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n902) );
  INV_X1 U676 ( .A(G1991), .ZN(n860) );
  NOR2_X1 U677 ( .A1(n902), .A2(n860), .ZN(n617) );
  XOR2_X1 U678 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n609) );
  NAND2_X1 U679 ( .A1(G105), .A2(n892), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G117), .A2(n888), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G129), .A2(n889), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n591), .A2(G141), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n884) );
  AND2_X1 U687 ( .A1(n884), .A2(G1996), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n940) );
  INV_X1 U689 ( .A(n940), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n618), .A2(n757), .ZN(n745) );
  NAND2_X1 U691 ( .A1(n752), .A2(n745), .ZN(n741) );
  XNOR2_X1 U692 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n674) );
  XNOR2_X1 U693 ( .A(KEYINPUT89), .B(n619), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n646) );
  INV_X1 U695 ( .A(n646), .ZN(n675) );
  INV_X1 U696 ( .A(G2072), .ZN(n955) );
  NOR2_X1 U697 ( .A1(n659), .A2(n955), .ZN(n623) );
  XNOR2_X1 U698 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n659), .A2(G1956), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT93), .B(n626), .ZN(n668) );
  NAND2_X1 U703 ( .A1(G53), .A2(n801), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G65), .A2(n802), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G91), .A2(n805), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G78), .A2(n806), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n980) );
  NOR2_X1 U710 ( .A1(n668), .A2(n980), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(n672) );
  NAND2_X1 U712 ( .A1(G1996), .A2(n675), .ZN(n635) );
  XNOR2_X1 U713 ( .A(KEYINPUT26), .B(n635), .ZN(n650) );
  NAND2_X1 U714 ( .A1(G56), .A2(n802), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT14), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n805), .A2(G81), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(KEYINPUT12), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G68), .A2(n806), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U720 ( .A(KEYINPUT13), .B(n640), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n643), .B(KEYINPUT71), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G43), .A2(n801), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n990) );
  NAND2_X1 U724 ( .A1(n646), .A2(G1341), .ZN(n647) );
  XOR2_X1 U725 ( .A(KEYINPUT94), .B(n647), .Z(n648) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n664) );
  NAND2_X1 U727 ( .A1(G92), .A2(n805), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G79), .A2(n806), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G54), .A2(n801), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G66), .A2(n802), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U734 ( .A(n657), .B(KEYINPUT15), .Z(n985) );
  INV_X1 U735 ( .A(n985), .ZN(n786) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT95), .ZN(n663) );
  NAND2_X1 U737 ( .A1(G1348), .A2(n646), .ZN(n661) );
  NAND2_X1 U738 ( .A1(G2067), .A2(n677), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n664), .A2(n786), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(KEYINPUT96), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n668), .A2(n980), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n674), .B(n673), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n675), .A2(G1961), .ZN(n676) );
  XOR2_X1 U749 ( .A(KEYINPUT90), .B(n676), .Z(n679) );
  XNOR2_X1 U750 ( .A(G2078), .B(KEYINPUT25), .ZN(n950) );
  NAND2_X1 U751 ( .A1(n677), .A2(n950), .ZN(n678) );
  NAND2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n687), .A2(G171), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n681), .A2(n680), .ZN(n704) );
  XNOR2_X1 U755 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n691) );
  NAND2_X1 U756 ( .A1(G8), .A2(n646), .ZN(n731) );
  NOR2_X1 U757 ( .A1(G1966), .A2(n731), .ZN(n706) );
  NOR2_X1 U758 ( .A1(G2084), .A2(n646), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G8), .A2(n682), .ZN(n683) );
  XNOR2_X1 U761 ( .A(KEYINPUT30), .B(n683), .ZN(n684) );
  XNOR2_X1 U762 ( .A(n684), .B(KEYINPUT98), .ZN(n685) );
  NOR2_X1 U763 ( .A1(G168), .A2(n685), .ZN(n686) );
  XNOR2_X1 U764 ( .A(n686), .B(KEYINPUT99), .ZN(n689) );
  OR2_X1 U765 ( .A1(n687), .A2(G171), .ZN(n688) );
  NAND2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U767 ( .A(n691), .B(n690), .ZN(n703) );
  INV_X1 U768 ( .A(G8), .ZN(n696) );
  NOR2_X1 U769 ( .A1(G2090), .A2(n646), .ZN(n693) );
  NOR2_X1 U770 ( .A1(G1971), .A2(n731), .ZN(n692) );
  NOR2_X1 U771 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U772 ( .A1(n694), .A2(G303), .ZN(n695) );
  OR2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n698) );
  AND2_X1 U774 ( .A1(n703), .A2(n698), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n704), .A2(n697), .ZN(n701) );
  INV_X1 U776 ( .A(n698), .ZN(n699) );
  OR2_X1 U777 ( .A1(n699), .A2(G286), .ZN(n700) );
  NAND2_X1 U778 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U779 ( .A(n702), .B(KEYINPUT32), .ZN(n711) );
  AND2_X1 U780 ( .A1(n704), .A2(n703), .ZN(n709) );
  AND2_X1 U781 ( .A1(G8), .A2(n705), .ZN(n707) );
  OR2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n727) );
  NOR2_X1 U784 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U785 ( .A1(G1971), .A2(G303), .ZN(n712) );
  XOR2_X1 U786 ( .A(n712), .B(KEYINPUT101), .Z(n713) );
  NOR2_X1 U787 ( .A1(n976), .A2(n713), .ZN(n714) );
  NAND2_X1 U788 ( .A1(n727), .A2(n714), .ZN(n715) );
  XNOR2_X1 U789 ( .A(n715), .B(KEYINPUT102), .ZN(n721) );
  NAND2_X1 U790 ( .A1(G1976), .A2(G288), .ZN(n978) );
  INV_X1 U791 ( .A(n978), .ZN(n716) );
  NOR2_X1 U792 ( .A1(n731), .A2(n716), .ZN(n718) );
  NAND2_X1 U793 ( .A1(n976), .A2(KEYINPUT33), .ZN(n717) );
  OR2_X1 U794 ( .A1(n717), .A2(n731), .ZN(n722) );
  AND2_X1 U795 ( .A1(n718), .A2(n722), .ZN(n719) );
  XOR2_X1 U796 ( .A(G1981), .B(G305), .Z(n973) );
  AND2_X1 U797 ( .A1(n719), .A2(n973), .ZN(n720) );
  AND2_X1 U798 ( .A1(n721), .A2(n720), .ZN(n737) );
  INV_X1 U799 ( .A(n973), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n722), .A2(KEYINPUT33), .ZN(n723) );
  OR2_X1 U801 ( .A1(n724), .A2(n723), .ZN(n735) );
  NOR2_X1 U802 ( .A1(G2090), .A2(G303), .ZN(n725) );
  NAND2_X1 U803 ( .A1(G8), .A2(n725), .ZN(n726) );
  NAND2_X1 U804 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U805 ( .A1(n728), .A2(n731), .ZN(n733) );
  NOR2_X1 U806 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XOR2_X1 U807 ( .A(n729), .B(KEYINPUT24), .Z(n730) );
  OR2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n744) );
  XOR2_X1 U812 ( .A(G1986), .B(G290), .Z(n742) );
  XNOR2_X1 U813 ( .A(KEYINPUT85), .B(n742), .ZN(n996) );
  NAND2_X1 U814 ( .A1(n996), .A2(n757), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n760) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n884), .ZN(n935) );
  INV_X1 U817 ( .A(n745), .ZN(n749) );
  AND2_X1 U818 ( .A1(n860), .A2(n902), .ZN(n941) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n746) );
  XNOR2_X1 U820 ( .A(KEYINPUT104), .B(n746), .ZN(n747) );
  NOR2_X1 U821 ( .A1(n941), .A2(n747), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n935), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U826 ( .A(KEYINPUT105), .B(n754), .Z(n756) );
  NAND2_X1 U827 ( .A1(n903), .A2(n755), .ZN(n927) );
  NAND2_X1 U828 ( .A1(n756), .A2(n927), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U831 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U832 ( .A(G2435), .B(G2446), .Z(n763) );
  XNOR2_X1 U833 ( .A(KEYINPUT106), .B(G2451), .ZN(n762) );
  XNOR2_X1 U834 ( .A(n763), .B(n762), .ZN(n767) );
  XOR2_X1 U835 ( .A(G2438), .B(KEYINPUT108), .Z(n765) );
  XNOR2_X1 U836 ( .A(KEYINPUT107), .B(G2454), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n765), .B(n764), .ZN(n766) );
  XOR2_X1 U838 ( .A(n767), .B(n766), .Z(n769) );
  XNOR2_X1 U839 ( .A(G2443), .B(G2427), .ZN(n768) );
  XNOR2_X1 U840 ( .A(n769), .B(n768), .ZN(n772) );
  XOR2_X1 U841 ( .A(G1341), .B(G1348), .Z(n770) );
  XNOR2_X1 U842 ( .A(G2430), .B(n770), .ZN(n771) );
  XOR2_X1 U843 ( .A(n772), .B(n771), .Z(n773) );
  AND2_X1 U844 ( .A1(G14), .A2(n773), .ZN(G401) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U846 ( .A1(G123), .A2(n889), .ZN(n774) );
  XNOR2_X1 U847 ( .A(n774), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U848 ( .A1(G111), .A2(n888), .ZN(n776) );
  NAND2_X1 U849 ( .A1(G135), .A2(n591), .ZN(n775) );
  NAND2_X1 U850 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U851 ( .A1(G99), .A2(n892), .ZN(n777) );
  XNOR2_X1 U852 ( .A(KEYINPUT75), .B(n777), .ZN(n778) );
  NOR2_X1 U853 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U854 ( .A1(n781), .A2(n780), .ZN(n931) );
  XNOR2_X1 U855 ( .A(G2096), .B(n931), .ZN(n782) );
  OR2_X1 U856 ( .A1(G2100), .A2(n782), .ZN(G156) );
  INV_X1 U857 ( .A(G132), .ZN(G219) );
  INV_X1 U858 ( .A(G82), .ZN(G220) );
  INV_X1 U859 ( .A(G120), .ZN(G236) );
  INV_X1 U860 ( .A(G69), .ZN(G235) );
  XOR2_X1 U861 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n785) );
  NAND2_X1 U862 ( .A1(G7), .A2(G661), .ZN(n783) );
  XOR2_X1 U863 ( .A(n783), .B(KEYINPUT10), .Z(n840) );
  NAND2_X1 U864 ( .A1(G567), .A2(n840), .ZN(n784) );
  XNOR2_X1 U865 ( .A(n785), .B(n784), .ZN(G234) );
  INV_X1 U866 ( .A(G860), .ZN(n792) );
  OR2_X1 U867 ( .A1(n990), .A2(n792), .ZN(G153) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n788) );
  INV_X1 U869 ( .A(G868), .ZN(n822) );
  NAND2_X1 U870 ( .A1(n786), .A2(n822), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n788), .A2(n787), .ZN(G284) );
  NAND2_X1 U872 ( .A1(n980), .A2(n822), .ZN(n789) );
  XNOR2_X1 U873 ( .A(n789), .B(KEYINPUT73), .ZN(n791) );
  NOR2_X1 U874 ( .A1(n822), .A2(G286), .ZN(n790) );
  NOR2_X1 U875 ( .A1(n791), .A2(n790), .ZN(G297) );
  NAND2_X1 U876 ( .A1(n792), .A2(G559), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n793), .A2(n985), .ZN(n794) );
  XNOR2_X1 U878 ( .A(n794), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n990), .ZN(n795) );
  XNOR2_X1 U880 ( .A(KEYINPUT74), .B(n795), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G868), .A2(n985), .ZN(n796) );
  NOR2_X1 U882 ( .A1(G559), .A2(n796), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(G282) );
  XNOR2_X1 U884 ( .A(n990), .B(KEYINPUT76), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n985), .A2(G559), .ZN(n799) );
  XNOR2_X1 U886 ( .A(n800), .B(n799), .ZN(n819) );
  NOR2_X1 U887 ( .A1(G860), .A2(n819), .ZN(n812) );
  NAND2_X1 U888 ( .A1(G55), .A2(n801), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G67), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n811) );
  NAND2_X1 U891 ( .A1(G93), .A2(n805), .ZN(n808) );
  NAND2_X1 U892 ( .A1(G80), .A2(n806), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U894 ( .A(KEYINPUT77), .B(n809), .Z(n810) );
  OR2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n821) );
  XOR2_X1 U896 ( .A(n812), .B(n821), .Z(G145) );
  INV_X1 U897 ( .A(n980), .ZN(G299) );
  XOR2_X1 U898 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n814) );
  XOR2_X1 U899 ( .A(G299), .B(G288), .Z(n813) );
  XNOR2_X1 U900 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n815), .B(n821), .ZN(n817) );
  XOR2_X1 U902 ( .A(G290), .B(G303), .Z(n816) );
  XNOR2_X1 U903 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U904 ( .A(n818), .B(G305), .ZN(n908) );
  XNOR2_X1 U905 ( .A(n819), .B(n908), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n820), .A2(G868), .ZN(n824) );
  NAND2_X1 U907 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U908 ( .A1(n824), .A2(n823), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2084), .A2(G2078), .ZN(n827) );
  XNOR2_X1 U910 ( .A(KEYINPUT81), .B(KEYINPUT20), .ZN(n825) );
  XNOR2_X1 U911 ( .A(n825), .B(KEYINPUT82), .ZN(n826) );
  XNOR2_X1 U912 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U913 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G235), .A2(G236), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT83), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G237), .A2(n832), .ZN(n833) );
  NAND2_X1 U921 ( .A1(G108), .A2(n833), .ZN(n844) );
  NAND2_X1 U922 ( .A1(n844), .A2(G567), .ZN(n838) );
  NOR2_X1 U923 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U924 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U925 ( .A1(G218), .A2(n835), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G96), .A2(n836), .ZN(n845) );
  NAND2_X1 U927 ( .A1(n845), .A2(G2106), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(n919) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n839) );
  NOR2_X1 U930 ( .A1(n919), .A2(n839), .ZN(n843) );
  NAND2_X1 U931 ( .A1(n843), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n840), .ZN(G217) );
  INV_X1 U933 ( .A(n840), .ZN(G223) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U935 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U939 ( .A(G108), .ZN(G238) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2084), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n846), .B(G2096), .ZN(n856) );
  XOR2_X1 U945 ( .A(G2678), .B(KEYINPUT110), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2100), .B(KEYINPUT109), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XOR2_X1 U949 ( .A(G2078), .B(n955), .Z(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n859), .B(G2474), .Z(n862) );
  XOR2_X1 U959 ( .A(G1996), .B(n860), .Z(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(KEYINPUT41), .B(G1981), .Z(n864) );
  XNOR2_X1 U962 ( .A(G1961), .B(G1956), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G124), .A2(n889), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n888), .A2(G112), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G136), .A2(n591), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G100), .A2(n892), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G139), .A2(n591), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G103), .A2(n892), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G115), .A2(n888), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G127), .A2(n889), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n920) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n882) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(n883), .B(G162), .Z(n886) );
  XOR2_X1 U985 ( .A(G160), .B(n884), .Z(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U987 ( .A(G164), .B(n887), .ZN(n900) );
  NAND2_X1 U988 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U991 ( .A1(G142), .A2(n591), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G106), .A2(n892), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(n895), .B(KEYINPUT45), .Z(n896) );
  NOR2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n898), .B(n931), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n920), .B(n901), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1002 ( .A(G286), .B(G171), .Z(n907) );
  XOR2_X1 U1003 ( .A(n907), .B(n985), .Z(n910) );
  XOR2_X1 U1004 ( .A(n990), .B(n908), .Z(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n912), .Z(n915) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n919), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT114), .B(n913), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(n916), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n919), .ZN(G319) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n948) );
  XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n926) );
  XNOR2_X1 U1019 ( .A(G164), .B(G2078), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n920), .B(KEYINPUT117), .ZN(n921) );
  XOR2_X1 U1021 ( .A(n921), .B(G2072), .Z(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT119), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n926), .B(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n944) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT116), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT51), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  XOR2_X1 U1038 ( .A(KEYINPUT120), .B(n946), .Z(n947) );
  NAND2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1040 ( .A1(n949), .A2(G29), .ZN(n1002) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1042 ( .A(n950), .B(G27), .Z(n952) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT122), .B(n953), .ZN(n960) );
  XOR2_X1 U1046 ( .A(G25), .B(G1991), .Z(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(n955), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G33), .B(n956), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(n969), .Z(n971) );
  INV_X1 U1060 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n972), .ZN(n1000) );
  XOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .Z(n998) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(KEYINPUT57), .ZN(n994) );
  INV_X1 U1067 ( .A(n976), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n979), .B(KEYINPUT123), .ZN(n989) );
  XOR2_X1 U1070 ( .A(G301), .B(G1961), .Z(n984) );
  XOR2_X1 U1071 ( .A(n980), .B(G1956), .Z(n982) );
  XOR2_X1 U1072 ( .A(G166), .B(G1971), .Z(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1075 ( .A(G1348), .B(n985), .Z(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1082 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1083 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1084 ( .A1(n1002), .A2(n1001), .ZN(n1029) );
  XOR2_X1 U1085 ( .A(G1961), .B(KEYINPUT124), .Z(n1003) );
  XNOR2_X1 U1086 ( .A(G5), .B(n1003), .ZN(n1023) );
  XOR2_X1 U1087 ( .A(G1966), .B(G21), .Z(n1014) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n1004), .B(G4), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G19), .B(G1341), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(G1981), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(G6), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(n1024), .B(KEYINPUT61), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(n1025), .B(KEYINPUT126), .ZN(n1026) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1026), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1027), .Z(n1028) );
  NOR2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1030), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

