//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n188));
  INV_X1    g002(.A(G122), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT92), .A3(G122), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT14), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n196), .A3(new_n192), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT78), .A2(G107), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT78), .A2(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n193), .A2(new_n203), .A3(new_n195), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n208), .A3(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n199), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT13), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n216), .A3(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n212), .A3(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n206), .A2(new_n208), .A3(new_n216), .A4(G134), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n203), .B1(new_n193), .B2(new_n195), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n219), .C1(new_n204), .C2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT9), .B(G234), .ZN(new_n222));
  INV_X1    g036(.A(G217), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n222), .A2(new_n223), .A3(G953), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n215), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n215), .B2(new_n221), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n187), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT93), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G478), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT15), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT93), .B(new_n187), .C1(new_n225), .C2(new_n226), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT94), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n227), .A2(new_n231), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n234), .B1(new_n233), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(G234), .A2(G237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(G902), .A3(G953), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT21), .B(G898), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n243), .A2(G952), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n242), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G113), .B(G122), .ZN(new_n247));
  INV_X1    g061(.A(G104), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n243), .A3(G214), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n205), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT18), .A2(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT18), .A2(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G140), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G140), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT89), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(KEYINPUT72), .A3(G125), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n264), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n260), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n270), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(G146), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n274), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT90), .A3(new_n260), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n266), .A2(KEYINPUT16), .A3(new_n268), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT16), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n262), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n271), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n255), .A2(G131), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n252), .A2(new_n290), .A3(new_n254), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n278), .A2(KEYINPUT19), .A3(new_n279), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(KEYINPUT19), .B2(new_n273), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n294), .B2(G146), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n249), .B1(new_n284), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n297), .A3(new_n291), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n255), .A2(KEYINPUT17), .A3(G131), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n285), .A2(new_n271), .A3(new_n287), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n288), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n285), .A2(new_n287), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT73), .A3(G146), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n300), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n275), .A2(new_n276), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT90), .B1(new_n282), .B2(new_n260), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n308), .B(new_n249), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT91), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n284), .A2(new_n313), .A3(new_n249), .A4(new_n308), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n296), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G475), .A2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT20), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n296), .ZN(new_n319));
  INV_X1    g133(.A(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n305), .A2(G146), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n302), .A3(new_n301), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n306), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n277), .A2(new_n283), .B1(new_n323), .B2(new_n300), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n313), .B1(new_n324), .B2(new_n249), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n319), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n316), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n320), .A2(new_n325), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n324), .A2(new_n249), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n187), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n318), .A2(new_n328), .B1(new_n331), .B2(G475), .ZN(new_n332));
  OAI21_X1  g146(.A(G221), .B1(new_n222), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n243), .A2(G227), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT77), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G143), .B(G146), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n271), .A2(G143), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n207), .B1(new_n343), .B2(KEYINPUT1), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(KEYINPUT78), .A2(G107), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G104), .A4(new_n200), .ZN(new_n348));
  INV_X1    g162(.A(G107), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n349), .B2(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(G104), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G101), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(G104), .B1(new_n346), .B2(new_n200), .ZN(new_n355));
  INV_X1    g169(.A(new_n351), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n248), .B1(new_n201), .B2(new_n202), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n353), .B1(new_n360), .B2(new_n351), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT65), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n205), .B2(G146), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n271), .A2(KEYINPUT65), .A3(G143), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n205), .A2(G146), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n205), .A2(G146), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n369));
  OAI21_X1  g183(.A(G128), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n342), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n358), .B1(new_n362), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n210), .A2(G137), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n210), .A2(G137), .ZN(new_n379));
  INV_X1    g193(.A(G137), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G134), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n381), .B2(new_n374), .ZN(new_n382));
  OAI21_X1  g196(.A(G131), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(G134), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n375), .B2(new_n376), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n374), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n290), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n373), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT12), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n373), .A2(KEYINPUT12), .A3(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT79), .B1(new_n359), .B2(new_n361), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n357), .A2(new_n354), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n395), .A2(KEYINPUT10), .A3(new_n372), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n348), .A2(new_n352), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n354), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT0), .A2(G128), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT0), .A2(G128), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n367), .A2(new_n404), .B1(new_n402), .B2(new_n340), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n406), .A3(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n389), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n358), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n398), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n339), .B1(new_n394), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n412), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n407), .A2(new_n405), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n415), .A2(new_n401), .B1(new_n410), .B2(new_n358), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n409), .B1(new_n416), .B2(new_n398), .ZN(new_n417));
  INV_X1    g231(.A(new_n339), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n335), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n393), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT12), .B1(new_n373), .B2(new_n389), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n412), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n418), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n412), .A2(new_n339), .ZN(new_n425));
  INV_X1    g239(.A(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(KEYINPUT80), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(G469), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n187), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n394), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n418), .B1(new_n414), .B2(new_n417), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n334), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n246), .A2(new_n332), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n443));
  AOI221_X4 g257(.A(G125), .B1(new_n340), .B2(new_n341), .C1(new_n367), .C2(new_n370), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n367), .A2(new_n404), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n340), .A2(new_n402), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n263), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n443), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n371), .A2(new_n263), .A3(new_n342), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n263), .B2(new_n405), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n443), .ZN(new_n453));
  INV_X1    g267(.A(G119), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G116), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(G113), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n191), .A2(G119), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n456), .B2(new_n457), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT2), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT67), .B1(new_n467), .B2(new_n457), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT2), .A3(G113), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n468), .A2(new_n470), .B1(new_n467), .B2(new_n457), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n462), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n362), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT8), .Z(new_n476));
  AOI22_X1  g290(.A1(new_n463), .A2(new_n458), .B1(new_n471), .B2(new_n462), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n357), .A2(new_n354), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n450), .A2(new_n453), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n445), .A2(new_n446), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT83), .B1(new_n482), .B2(G125), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n452), .B2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g298(.A(new_n443), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT86), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT83), .B1(new_n444), .B2(new_n447), .ZN(new_n487));
  INV_X1    g301(.A(new_n483), .ZN(new_n488));
  AND4_X1   g302(.A1(KEYINPUT86), .A2(new_n487), .A3(new_n488), .A4(new_n485), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n480), .B(new_n481), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n395), .A2(new_n477), .A3(new_n397), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n468), .A2(new_n470), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n467), .A2(new_n457), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n461), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n472), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n401), .A2(new_n496), .A3(new_n407), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n497), .A3(new_n475), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n487), .A2(new_n488), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n443), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n484), .A2(KEYINPUT86), .A3(new_n485), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n481), .B1(new_n504), .B2(new_n480), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n491), .A2(new_n497), .ZN(new_n507));
  INV_X1    g321(.A(new_n475), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT82), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n498), .A2(new_n510), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n484), .B(new_n441), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n187), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n439), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n480), .B1(new_n486), .B2(new_n489), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n498), .A3(new_n490), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n513), .A2(new_n512), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n515), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n525), .A3(new_n438), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G214), .B1(G237), .B2(G902), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT81), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n520), .A2(new_n525), .A3(new_n438), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n527), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n437), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n378), .A2(new_n382), .A3(G131), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n290), .B1(new_n385), .B2(new_n387), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n405), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G131), .B1(new_n376), .B2(new_n384), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT65), .B1(new_n271), .B2(G143), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n271), .A2(G143), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n344), .B1(new_n542), .B2(new_n365), .ZN(new_n543));
  INV_X1    g357(.A(new_n342), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n388), .B(new_n539), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT30), .B1(new_n546), .B2(KEYINPUT64), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT64), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  AOI211_X1 g363(.A(new_n548), .B(new_n549), .C1(new_n538), .C2(new_n545), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n496), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT26), .B(G101), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n253), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n471), .B(new_n461), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n538), .A2(new_n558), .A3(new_n545), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n546), .A2(new_n496), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT69), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n556), .B(new_n563), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT31), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n551), .A2(KEYINPUT31), .A3(new_n557), .A4(new_n559), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n187), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n572), .A2(new_n187), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n571), .A4(new_n570), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n538), .A2(new_n558), .A3(new_n545), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n558), .B1(new_n538), .B2(new_n545), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT28), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT69), .A3(new_n566), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n556), .B1(new_n581), .B2(new_n563), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n582), .B2(KEYINPUT29), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n557), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n546), .A2(KEYINPUT64), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n549), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n546), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n558), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n556), .B1(new_n589), .B2(new_n578), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n574), .A2(new_n577), .B1(G472), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n223), .B1(G234), .B2(new_n187), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n454), .B2(G128), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n454), .A2(G128), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT70), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n598), .A2(new_n599), .A3(new_n603), .A4(new_n600), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(G110), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n605), .A2(KEYINPUT71), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n207), .A2(G119), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n600), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT24), .B(G110), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n605), .B2(KEYINPUT71), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n322), .A2(new_n606), .A3(new_n306), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(G110), .B2(new_n601), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n321), .A2(new_n613), .A3(new_n281), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n281), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT74), .B1(new_n617), .B2(new_n288), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT75), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT22), .B(G137), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n612), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n612), .B2(new_n619), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n187), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(KEYINPUT25), .B(new_n187), .C1(new_n624), .C2(new_n625), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n596), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n625), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n595), .A2(G902), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT76), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n594), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n535), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  NAND2_X1  g453(.A1(new_n328), .A2(new_n318), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n330), .B1(new_n312), .B2(new_n314), .ZN(new_n641));
  OAI21_X1  g455(.A(G475), .B1(new_n641), .B2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n229), .A2(new_n232), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(G478), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n225), .A2(new_n226), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT33), .B1(new_n226), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n230), .A2(G902), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n644), .A2(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n245), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n429), .A2(new_n435), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n635), .A3(new_n333), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n571), .B1(new_n575), .B2(new_n570), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n560), .A2(new_n568), .A3(new_n569), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n572), .A2(new_n187), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n659), .A2(G472), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT95), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT95), .A3(new_n573), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n657), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n529), .B1(new_n517), .B2(new_n526), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n655), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G104), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(new_n238), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n643), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n245), .B(KEYINPUT99), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NAND2_X1  g492(.A1(new_n628), .A2(new_n629), .ZN(new_n679));
  INV_X1    g493(.A(new_n633), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n612), .A2(new_n619), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n623), .A2(KEYINPUT36), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n679), .A2(new_n595), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n663), .B2(new_n665), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n535), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n574), .A2(new_n577), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n593), .A2(G472), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n244), .A2(new_n239), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT100), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(G900), .B2(new_n240), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n642), .A2(new_n640), .A3(new_n238), .A4(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n695), .A3(new_n436), .A4(new_n667), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  INV_X1    g511(.A(new_n684), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n694), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n436), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n529), .B(new_n698), .C1(new_n700), .C2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n551), .A2(new_n559), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n557), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n564), .A2(new_n556), .A3(new_n559), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n187), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n332), .A2(new_n672), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n701), .A2(new_n708), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n527), .A2(new_n533), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT38), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NAND2_X1  g529(.A1(new_n689), .A2(new_n690), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n436), .A3(new_n667), .A4(new_n698), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n643), .A2(new_n653), .A3(new_n694), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT101), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n656), .A2(new_n333), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n594), .A2(new_n720), .A3(new_n684), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  INV_X1    g536(.A(new_n694), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n652), .B(new_n723), .C1(new_n640), .C2(new_n642), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n722), .A3(new_n667), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  NAND2_X1  g541(.A1(new_n432), .A2(new_n433), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n187), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n434), .A2(new_n430), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n333), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n655), .A2(new_n637), .A3(new_n667), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n637), .A2(new_n675), .A3(new_n673), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AOI21_X1  g552(.A(new_n438), .B1(new_n520), .B2(new_n525), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n530), .B1(new_n531), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n732), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n691), .A3(new_n332), .A4(new_n246), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  AND4_X1   g557(.A1(new_n333), .A2(new_n730), .A3(new_n731), .A4(new_n674), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n643), .A2(new_n744), .A3(new_n667), .A4(new_n238), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n679), .A2(new_n595), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT102), .ZN(new_n747));
  INV_X1    g561(.A(new_n634), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT102), .B1(new_n630), .B2(new_n634), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n661), .A2(new_n658), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n745), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT104), .B(G122), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G24));
  AOI21_X1  g572(.A(KEYINPUT105), .B1(new_n753), .B2(new_n698), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n664), .A2(new_n573), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n760), .A2(new_n761), .A3(new_n684), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n724), .B(new_n741), .C1(new_n759), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  AOI21_X1  g578(.A(new_n529), .B1(new_n527), .B2(new_n533), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n413), .A2(new_n419), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(G469), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n413), .A2(new_n419), .A3(KEYINPUT106), .A4(new_n430), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n334), .B1(new_n771), .B2(new_n435), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n765), .B2(new_n772), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n637), .B(new_n724), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT108), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n712), .A2(new_n772), .A3(new_n530), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT107), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n653), .A4(new_n694), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n749), .A2(new_n750), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT109), .B1(new_n786), .B2(new_n594), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n716), .A2(new_n788), .A3(new_n751), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT110), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n784), .A2(new_n790), .A3(KEYINPUT110), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n778), .B(new_n780), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G131), .ZN(G33));
  OAI211_X1 g608(.A(new_n637), .B(new_n695), .C1(new_n773), .C2(new_n774), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT111), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n784), .A2(new_n797), .A3(new_n637), .A4(new_n695), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  INV_X1    g614(.A(new_n765), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(G469), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n420), .B2(new_n428), .ZN(new_n804));
  OAI22_X1  g618(.A1(new_n803), .A2(new_n804), .B1(new_n430), .B2(new_n187), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n805), .A2(new_n806), .B1(new_n430), .B2(new_n434), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n333), .A3(new_n699), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n332), .A2(new_n653), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT43), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(KEYINPUT112), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n332), .A2(new_n653), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n663), .A2(new_n665), .A3(new_n698), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n801), .B(new_n809), .C1(new_n810), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(KEYINPUT44), .A3(new_n817), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n333), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(KEYINPUT47), .A3(new_n333), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n718), .A2(new_n716), .A3(new_n635), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n765), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND3_X1  g644(.A1(new_n751), .A2(new_n530), .A3(new_n333), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n730), .A2(new_n731), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT49), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n811), .A3(new_n708), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n713), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n754), .A2(new_n755), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n693), .B1(new_n813), .B2(new_n815), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n713), .A2(new_n529), .A3(new_n733), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n801), .A2(new_n732), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n759), .A2(new_n762), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n708), .A2(new_n636), .A3(new_n692), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n332), .A2(new_n652), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n844), .A2(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n825), .B(new_n826), .C1(new_n333), .C2(new_n833), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n837), .A2(new_n765), .A3(new_n838), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  INV_X1    g669(.A(new_n741), .ZN(new_n856));
  OAI221_X1 g670(.A(new_n244), .B1(new_n654), .B2(new_n847), .C1(new_n839), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n787), .A2(new_n789), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n838), .A2(new_n860), .A3(new_n843), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n842), .A2(new_n853), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n865));
  OAI221_X1 g679(.A(new_n863), .B1(new_n858), .B2(new_n857), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(new_n762), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n761), .B1(new_n760), .B2(new_n684), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n718), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n773), .B2(new_n774), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n233), .A2(new_n235), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n723), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n640), .A2(new_n642), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT114), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n721), .A3(new_n765), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n734), .A2(new_n737), .A3(new_n742), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n640), .A2(new_n642), .A3(new_n872), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n332), .B2(new_n652), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n666), .A2(new_n534), .A3(new_n674), .A4(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n437), .B(new_n534), .C1(new_n637), .C2(new_n685), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n756), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n877), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n763), .A2(new_n696), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n719), .B2(new_n725), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n740), .A2(new_n332), .A3(new_n672), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n698), .A2(new_n723), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n887), .A2(new_n708), .A3(new_n772), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT52), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n763), .A2(new_n696), .ZN(new_n891));
  AND4_X1   g705(.A1(KEYINPUT52), .A2(new_n726), .A3(new_n891), .A4(new_n889), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n799), .B(new_n884), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n780), .B1(new_n792), .B2(new_n791), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n779), .B1(new_n775), .B2(new_n776), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n867), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n884), .A2(new_n799), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n726), .A2(new_n891), .A3(new_n889), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n889), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(new_n793), .A3(KEYINPUT53), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n897), .A2(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n855), .B(new_n866), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n836), .B1(new_n910), .B2(new_n911), .ZN(G75));
  XNOR2_X1  g726(.A(new_n523), .B(new_n524), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n905), .A2(G210), .A3(G902), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n243), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n915), .A2(KEYINPUT56), .A3(new_n914), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G51));
  XNOR2_X1  g735(.A(new_n431), .B(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n909), .A2(new_n907), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n728), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n908), .A2(new_n187), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n803), .A2(new_n804), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n924), .B2(new_n927), .ZN(G54));
  AND2_X1   g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n925), .A2(new_n326), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n326), .B1(new_n925), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n917), .ZN(G60));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT59), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n909), .A2(new_n907), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n650), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n917), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n909), .A2(new_n650), .A3(new_n907), .A4(new_n934), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n223), .A2(new_n187), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n905), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n631), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT119), .B1(new_n945), .B2(new_n918), .ZN(new_n946));
  INV_X1    g760(.A(new_n943), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n897), .B2(new_n904), .ZN(new_n948));
  INV_X1    g762(.A(new_n631), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT119), .B(new_n918), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n905), .A2(new_n683), .A3(new_n943), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n940), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n918), .B1(new_n948), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n940), .B1(new_n948), .B2(new_n683), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n945), .A2(new_n958), .A3(KEYINPUT120), .A4(new_n918), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n953), .A2(new_n960), .ZN(G66));
  NOR2_X1   g775(.A1(new_n883), .A2(new_n878), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(G953), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT121), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n242), .B2(new_n440), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n514), .B1(G898), .B2(new_n243), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  AND2_X1   g782(.A1(new_n821), .A2(new_n829), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n714), .A2(new_n886), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n972));
  INV_X1    g786(.A(new_n700), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n637), .A2(new_n880), .A3(new_n973), .A4(new_n765), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n243), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n547), .A2(new_n550), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n294), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n243), .A2(G900), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT123), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n860), .A2(new_n887), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n809), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n985), .A2(new_n886), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n969), .A3(new_n793), .A4(new_n799), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n987), .B2(new_n243), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n979), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT122), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n989), .B(new_n992), .ZN(G72));
  XNOR2_X1  g807(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n571), .A2(new_n187), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n962), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n975), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g814(.A(KEYINPUT126), .B(new_n996), .C1(new_n975), .C2(new_n997), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n704), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n702), .A2(new_n557), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n905), .A2(new_n703), .A3(new_n996), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n996), .B1(new_n987), .B2(new_n997), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n917), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(G57));
endmodule


