//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n449, new_n451, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  NAND2_X1  g023(.A1(G94), .A2(G452), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT70), .Z(G261));
  AOI22_X1  g034(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT71), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(new_n461), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n481), .B1(new_n484), .B2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n462), .B2(new_n463), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n463), .C2(new_n462), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT72), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT72), .A2(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n505), .B2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n507), .A2(new_n508), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n515), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n503), .A2(new_n504), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(KEYINPUT73), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT73), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n506), .A2(new_n509), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n513), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G52), .Z(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G90), .B1(new_n514), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  INV_X1    g116(.A(G77), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n519), .A2(new_n541), .B1(new_n542), .B2(new_n502), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI221_X1 g120(.A(KEYINPUT74), .B1(new_n542), .B2(new_n502), .C1(new_n519), .C2(new_n541), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(new_n522), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n519), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n522), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n506), .A2(G81), .A3(new_n509), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n509), .A2(G43), .A3(new_n512), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(KEYINPUT78), .A2(G78), .A3(G543), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n526), .A2(G65), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n562), .B1(new_n567), .B2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  INV_X1    g144(.A(new_n566), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT78), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n503), .B2(new_n504), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n509), .A2(new_n512), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n509), .A2(new_n580), .A3(new_n512), .A4(new_n577), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n568), .A2(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n505), .A2(G651), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n509), .A2(new_n526), .A3(G91), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n506), .A2(new_n586), .A3(new_n509), .A4(G91), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n588), .ZN(G299));
  OAI21_X1  g164(.A(KEYINPUT80), .B1(new_n533), .B2(new_n537), .ZN(new_n590));
  INV_X1    g165(.A(new_n537), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n510), .A2(G89), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n526), .A2(new_n527), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n528), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G286));
  OAI21_X1  g175(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n509), .A2(G49), .A3(new_n512), .ZN(new_n602));
  INV_X1    g177(.A(G87), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n531), .C2(new_n603), .ZN(G288));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n519), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g182(.A(KEYINPUT81), .B(G61), .C1(new_n517), .C2(new_n518), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(new_n522), .B1(G48), .B2(new_n514), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n509), .A2(new_n526), .A3(G86), .A4(new_n583), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n506), .A2(KEYINPUT83), .A3(new_n509), .A4(G86), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n618), .A3(KEYINPUT84), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(KEYINPUT84), .B1(new_n613), .B2(new_n618), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(G305));
  NAND2_X1  g197(.A1(new_n510), .A2(G85), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n514), .A2(G47), .ZN(new_n624));
  NAND2_X1  g199(.A1(G72), .A2(G543), .ZN(new_n625));
  INV_X1    g200(.A(G60), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n519), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n522), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(G290));
  NAND2_X1  g204(.A1(G301), .A2(G868), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n631));
  INV_X1    g206(.A(G54), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n631), .A2(new_n562), .B1(new_n513), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n635));
  INV_X1    g210(.A(G92), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n531), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n630), .B1(G868), .B2(new_n638), .ZN(G321));
  XOR2_X1   g214(.A(G321), .B(KEYINPUT85), .Z(G284));
  NOR2_X1   g215(.A1(G299), .A2(G868), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n599), .ZN(G297));
  AOI21_X1  g217(.A(new_n641), .B1(G868), .B2(new_n599), .ZN(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n638), .B1(new_n644), .B2(G860), .ZN(G148));
  INV_X1    g220(.A(new_n638), .ZN(new_n646));
  OAI21_X1  g221(.A(KEYINPUT86), .B1(new_n646), .B2(G559), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G868), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n646), .A2(KEYINPUT86), .A3(G559), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n649), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n474), .A2(new_n468), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(G2100), .ZN(new_n658));
  OAI21_X1  g233(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n461), .A2(KEYINPUT87), .A3(G111), .ZN(new_n663));
  OAI21_X1  g238(.A(KEYINPUT87), .B1(new_n461), .B2(G111), .ZN(new_n664));
  NAND4_X1  g239(.A1(new_n661), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n484), .A2(G123), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n477), .B2(G135), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(G2096), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n657), .A2(G2100), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(G2096), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n658), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(G156));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2427), .B(G2438), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2430), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1341), .B(G1348), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n687), .A3(G14), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G401));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XOR2_X1   g266(.A(G2072), .B(G2078), .Z(new_n692));
  XNOR2_X1  g267(.A(G2084), .B(G2090), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT18), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(KEYINPUT17), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n696), .B(new_n693), .C1(new_n691), .C2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n693), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n691), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G2096), .B(G2100), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n695), .A2(new_n698), .A3(new_n700), .A4(new_n702), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(G227));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1971), .B(G1976), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT19), .ZN(new_n710));
  XOR2_X1   g285(.A(G1956), .B(G2474), .Z(new_n711));
  XOR2_X1   g286(.A(G1961), .B(G1966), .Z(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT20), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n712), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n710), .A2(new_n713), .A3(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G1981), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n714), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n717), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1981), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT90), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n720), .A2(new_n726), .A3(G1986), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n732), .B1(new_n729), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n708), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n729), .A2(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(new_n731), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(new_n739), .A3(new_n707), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(G229));
  INV_X1    g316(.A(KEYINPUT102), .ZN(new_n742));
  NAND2_X1  g317(.A1(G305), .A2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G6), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT32), .B(G1981), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n747), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n743), .A2(new_n749), .A3(new_n745), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n744), .A2(G22), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G303), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1971), .ZN(new_n753));
  MUX2_X1   g328(.A(G23), .B(G288), .S(G16), .Z(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT33), .B(G1976), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n748), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT34), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT34), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n748), .A2(new_n761), .A3(new_n750), .A4(new_n758), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G25), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n477), .A2(G131), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  INV_X1    g341(.A(G107), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G2105), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n484), .B2(G119), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n763), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT35), .B(G1991), .Z(new_n773));
  XOR2_X1   g348(.A(new_n772), .B(new_n773), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n744), .A2(G24), .ZN(new_n775));
  INV_X1    g350(.A(G290), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n744), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1986), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n760), .A2(new_n762), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(KEYINPUT36), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n760), .A2(new_n762), .A3(new_n782), .A4(new_n779), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n477), .A2(G140), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n786));
  INV_X1    g361(.A(G116), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G2105), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n484), .B2(G128), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n763), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n763), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT28), .Z(new_n792));
  OR3_X1    g367(.A1(new_n790), .A2(KEYINPUT91), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT91), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2067), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n793), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n744), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT23), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n763), .A2(G32), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n468), .A2(G105), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT26), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n805), .B(new_n807), .C1(G129), .C2(new_n484), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n477), .A2(G141), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT27), .B(G1996), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n744), .A2(G19), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n556), .B2(new_n744), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(G1341), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n763), .A2(G35), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n486), .B2(G29), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT29), .B(G2090), .Z(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n814), .A2(G1341), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n815), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n744), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n744), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G1961), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n763), .A2(G27), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G164), .B2(new_n763), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(G2078), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  AND2_X1   g406(.A1(KEYINPUT24), .A2(G34), .ZN(new_n832));
  NOR2_X1   g407(.A1(KEYINPUT24), .A2(G34), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n763), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT95), .Z(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G160), .B2(G29), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G2084), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n825), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n799), .A2(new_n803), .A3(new_n822), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n477), .A2(KEYINPUT92), .A3(G139), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n473), .A2(new_n476), .ZN(new_n843));
  INV_X1    g418(.A(G139), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT25), .Z(new_n847));
  NAND3_X1  g422(.A1(new_n841), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT93), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n461), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT94), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n848), .B2(KEYINPUT93), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G29), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n763), .A2(G33), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n442), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n840), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n744), .A2(G21), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G168), .B2(new_n744), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G1966), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT31), .B(G11), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT97), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT30), .B(G28), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(new_n763), .ZN(new_n866));
  AOI211_X1 g441(.A(new_n864), .B(new_n866), .C1(new_n668), .C2(G29), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n824), .A2(G1961), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n861), .A2(G1966), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT98), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n811), .A2(new_n812), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT96), .Z(new_n874));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n868), .A2(new_n875), .A3(new_n869), .A4(new_n870), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n744), .A2(G4), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n638), .B2(new_n744), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G1348), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n836), .A2(new_n880), .A3(G2084), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n836), .B2(G2084), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n818), .B2(new_n819), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AND4_X1   g459(.A1(new_n872), .A2(new_n874), .A3(new_n876), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n856), .A2(new_n442), .A3(new_n857), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n859), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n742), .B1(new_n784), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g464(.A(KEYINPUT102), .B(new_n887), .C1(new_n781), .C2(new_n783), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(G311));
  NAND2_X1  g466(.A1(new_n784), .A2(new_n888), .ZN(G150));
  NAND2_X1  g467(.A1(new_n638), .A2(G559), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT38), .Z(new_n894));
  NAND3_X1  g469(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n506), .A2(G93), .A3(new_n509), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n509), .A2(G55), .A3(new_n512), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n507), .A2(new_n508), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n895), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n894), .B(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT103), .B(G860), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT37), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(G145));
  XOR2_X1   g485(.A(new_n668), .B(G160), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n486), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n497), .A2(new_n499), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n488), .A2(new_n492), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g493(.A1(G164), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n484), .A2(G130), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n477), .A2(G142), .ZN(new_n923));
  OR3_X1    g498(.A1(new_n461), .A2(KEYINPUT106), .A3(G118), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n461), .B2(G118), .ZN(new_n925));
  OR2_X1    g500(.A1(G106), .A2(G2105), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n924), .A2(G2104), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n655), .B1(new_n765), .B2(new_n769), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n765), .A2(new_n655), .A3(new_n769), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n934), .B2(new_n930), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n920), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n785), .A2(new_n789), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n810), .B(new_n938), .Z(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n933), .A2(new_n935), .A3(new_n920), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n936), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n944), .A3(new_n854), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n854), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n913), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n912), .A4(new_n945), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g528(.A(new_n901), .B1(new_n648), .B2(new_n650), .ZN(new_n954));
  INV_X1    g529(.A(new_n650), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n556), .B(new_n900), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n647), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n646), .A2(G299), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n638), .A2(new_n588), .A3(new_n582), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n961), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT41), .B1(new_n960), .B2(new_n961), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n954), .A3(new_n957), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n959), .B1(new_n958), .B2(new_n962), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT110), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n969), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n967), .A4(new_n963), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n620), .A2(new_n621), .A3(new_n776), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n613), .A2(new_n618), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT84), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G290), .B1(new_n978), .B2(new_n619), .ZN(new_n979));
  XNOR2_X1  g554(.A(G303), .B(G288), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n975), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n776), .B1(new_n620), .B2(new_n621), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n619), .A3(G290), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n974), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n975), .B2(new_n979), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n980), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(KEYINPUT109), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n982), .B2(new_n985), .ZN(new_n993));
  AND4_X1   g568(.A1(new_n970), .A2(new_n973), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n970), .A2(new_n973), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(G868), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n900), .A2(new_n649), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(G295));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n997), .ZN(G331));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  AOI22_X1  g576(.A1(G89), .A2(new_n510), .B1(new_n596), .B2(new_n528), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n547), .A2(new_n540), .B1(new_n1002), .B2(new_n591), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(G171), .B2(new_n599), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n1004), .B2(new_n956), .ZN(new_n1005));
  AOI21_X1  g580(.A(G301), .B1(new_n590), .B2(new_n598), .ZN(new_n1006));
  NOR4_X1   g581(.A1(new_n1006), .A2(new_n901), .A3(new_n1003), .A4(KEYINPUT112), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n901), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n962), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n599), .A2(G171), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1003), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n956), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1009), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1008), .A2(new_n1010), .B1(new_n966), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G37), .B1(new_n990), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(KEYINPUT112), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1004), .A2(new_n1001), .A3(new_n956), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n1009), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n966), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(new_n989), .A3(new_n986), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1000), .B1(new_n1024), .B2(KEYINPUT43), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n951), .B1(new_n990), .B2(new_n1015), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT113), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n990), .A2(new_n1015), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n951), .C1(new_n990), .C2(new_n1015), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1031), .B2(KEYINPUT43), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1016), .A2(new_n1023), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n1031), .B2(KEYINPUT43), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n582), .B2(new_n588), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n579), .A2(new_n581), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n565), .A2(new_n566), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(KEYINPUT79), .C1(new_n519), .C2(new_n573), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n575), .A2(new_n1042), .A3(G651), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1038), .A2(new_n588), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n914), .B2(new_n915), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G40), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n466), .A2(new_n470), .A3(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1046), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G160), .A2(G40), .ZN(new_n1056));
  INV_X1    g631(.A(G1384), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n916), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(G1384), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n917), .A2(new_n919), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1045), .A2(new_n1055), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1039), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1044), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1064), .A2(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1069));
  INV_X1    g644(.A(new_n499), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n498), .B1(new_n474), .B2(new_n495), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1057), .B(new_n1053), .C1(new_n1072), .C2(new_n493), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1052), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1047), .A2(new_n797), .A3(new_n1052), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n646), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1065), .B1(new_n1068), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1045), .A2(new_n1055), .A3(new_n1064), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1068), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT122), .B(new_n1080), .C1(new_n1081), .C2(new_n1068), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n646), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n638), .A4(new_n1077), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1064), .A2(new_n1055), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1045), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1060), .A2(new_n1062), .A3(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1058), .B2(new_n1056), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1102), .B2(new_n556), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n895), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1092), .B(new_n1096), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1079), .B1(new_n1086), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1966), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1061), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(G164), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1061), .C1(new_n1072), .C2(new_n493), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT118), .B(new_n1052), .C1(new_n1047), .C2(KEYINPUT45), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1059), .B1(G164), .B2(G1384), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT118), .B1(new_n1115), .B2(new_n1052), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1069), .A2(new_n1073), .A3(new_n1118), .A4(new_n1052), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1056), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1122), .A2(KEYINPUT120), .A3(new_n1118), .A4(new_n1069), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1117), .A2(G168), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G8), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1126));
  AOI21_X1  g701(.A(G168), .B1(new_n1126), .B2(new_n1117), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT51), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1129), .A3(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(G2078), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1062), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n917), .A2(new_n919), .A3(new_n1057), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1059), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n1136), .B2(new_n1052), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n1056), .C1(new_n1135), .C2(new_n1059), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1060), .A2(new_n1062), .A3(new_n443), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1132), .ZN(new_n1142));
  INV_X1    g717(.A(G1961), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1074), .A2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(new_n1145), .A3(G301), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1116), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n1113), .A3(new_n1112), .A4(new_n1133), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G171), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1148), .A2(new_n1142), .A3(G301), .A4(new_n1144), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1155), .A2(KEYINPUT54), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1151), .A2(new_n1152), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1971), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1074), .A2(G2090), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1162), .B(G8), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G8), .ZN(new_n1166));
  INV_X1    g741(.A(G1971), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n917), .A2(new_n919), .A3(new_n1061), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1115), .A2(new_n1052), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1171));
  INV_X1    g746(.A(G2090), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1052), .A4(new_n1049), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1166), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1165), .B1(new_n1174), .B2(new_n1162), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT49), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n611), .A2(new_n608), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT81), .B1(new_n526), .B2(G61), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n522), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n514), .A2(G48), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n616), .A2(new_n617), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1181), .A2(G1981), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n725), .B1(new_n613), .B2(new_n614), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n614), .ZN(new_n1186));
  OAI21_X1  g761(.A(G1981), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1187), .B(KEYINPUT49), .C1(new_n976), .C2(G1981), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1166), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT52), .ZN(new_n1191));
  INV_X1    g766(.A(G1976), .ZN(new_n1192));
  OR2_X1    g767(.A1(G288), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT52), .B1(G288), .B2(new_n1192), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1158), .B1(new_n1175), .B2(new_n1198), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1173), .ZN(new_n1201));
  OAI21_X1  g776(.A(G8), .B1(new_n1201), .B2(new_n1163), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1161), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1203), .A2(new_n1159), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1200), .A2(new_n1205), .A3(KEYINPUT124), .A4(new_n1165), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1199), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1106), .A2(new_n1131), .A3(new_n1157), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1131), .A2(KEYINPUT62), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1128), .A2(new_n1210), .A3(new_n1130), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1150), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1199), .A2(new_n1206), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1209), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT117), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1165), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT116), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1190), .A2(new_n1217), .A3(new_n1197), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1217), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(G288), .A2(G1976), .ZN(new_n1221));
  AND2_X1   g796(.A1(new_n1190), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1189), .B1(new_n1222), .B2(new_n1183), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1215), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT63), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT121), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n599), .A2(G8), .ZN(new_n1227));
  AOI211_X1 g802(.A(new_n1226), .B(new_n1227), .C1(new_n1126), .C2(new_n1117), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1117), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1227), .ZN(new_n1230));
  AOI21_X1  g805(.A(KEYINPUT121), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1200), .A2(new_n1205), .A3(new_n1165), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1225), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1219), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1190), .A2(new_n1217), .A3(new_n1197), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1164), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1238), .A2(new_n1170), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1162), .B1(new_n1239), .B2(G8), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1165), .A2(KEYINPUT63), .ZN(new_n1241));
  NOR2_X1   g816(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g817(.A(new_n1237), .B(new_n1242), .C1(new_n1228), .C2(new_n1231), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1224), .B1(new_n1234), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g819(.A1(new_n1220), .A2(new_n1215), .A3(new_n1223), .ZN(new_n1245));
  NAND4_X1  g820(.A1(new_n1208), .A2(new_n1214), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NOR2_X1   g821(.A1(new_n1136), .A2(new_n1056), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n938), .A2(G2067), .ZN(new_n1248));
  NAND3_X1  g823(.A1(new_n785), .A2(new_n797), .A3(new_n789), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g825(.A(new_n1250), .B(KEYINPUT114), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n810), .B(new_n1098), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n771), .A2(new_n773), .ZN(new_n1253));
  OR2_X1    g828(.A1(new_n771), .A2(new_n773), .ZN(new_n1254));
  NAND4_X1  g829(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g830(.A(G290), .B(G1986), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1247), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1246), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g833(.A1(new_n1251), .A2(new_n809), .A3(new_n808), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1247), .A2(new_n1098), .ZN(new_n1260));
  OR2_X1    g835(.A1(new_n1260), .A2(KEYINPUT46), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1260), .A2(KEYINPUT46), .ZN(new_n1262));
  AOI22_X1  g837(.A1(new_n1247), .A2(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g838(.A(new_n1263), .B(KEYINPUT47), .Z(new_n1264));
  NAND3_X1  g839(.A1(new_n1247), .A2(new_n728), .A3(new_n776), .ZN(new_n1265));
  XNOR2_X1  g840(.A(new_n1265), .B(KEYINPUT125), .ZN(new_n1266));
  INV_X1    g841(.A(KEYINPUT48), .ZN(new_n1267));
  OR2_X1    g842(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g843(.A1(new_n1255), .A2(new_n1247), .ZN(new_n1269));
  NAND2_X1  g844(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1270));
  NAND3_X1  g845(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g846(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1272));
  OAI21_X1  g847(.A(new_n1249), .B1(new_n1272), .B2(new_n1253), .ZN(new_n1273));
  NAND2_X1  g848(.A1(new_n1273), .A2(new_n1247), .ZN(new_n1274));
  NAND3_X1  g849(.A1(new_n1264), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g850(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g851(.A1(new_n1258), .A2(new_n1276), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g852(.A1(new_n704), .A2(G319), .A3(new_n705), .ZN(new_n1279));
  XNOR2_X1  g853(.A(new_n1279), .B(KEYINPUT126), .ZN(new_n1280));
  AND3_X1   g854(.A1(new_n1280), .A2(KEYINPUT127), .A3(new_n688), .ZN(new_n1281));
  AOI21_X1  g855(.A(KEYINPUT127), .B1(new_n1280), .B2(new_n688), .ZN(new_n1282));
  NOR3_X1   g856(.A1(G229), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g857(.A1(new_n1283), .A2(new_n952), .ZN(new_n1284));
  NOR2_X1   g858(.A1(new_n1284), .A2(new_n1035), .ZN(G308));
  AND2_X1   g859(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1286));
  AOI21_X1  g860(.A(new_n1033), .B1(new_n1286), .B2(new_n1027), .ZN(new_n1287));
  OAI211_X1 g861(.A(new_n952), .B(new_n1283), .C1(new_n1287), .C2(new_n1034), .ZN(G225));
endmodule


