//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n464), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n472), .B1(new_n465), .B2(new_n466), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT68), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n473), .A2(new_n474), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n484), .B(new_n487), .C1(G136), .C2(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G138), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(new_n493), .A3(G138), .A4(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n472), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(G2104), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n498), .A2(new_n503), .B1(new_n485), .B2(G126), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(new_n511), .B1(new_n507), .B2(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n515), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(G51), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n521), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT71), .B(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n518), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n521), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n512), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n521), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n518), .A2(new_n559), .A3(G53), .ZN(new_n560));
  AND2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT6), .A2(G651), .ZN(new_n562));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n512), .A2(G91), .A3(new_n520), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n514), .ZN(G299));
  OR2_X1    g143(.A1(new_n515), .A2(new_n523), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n512), .A2(G87), .A3(new_n520), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n518), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n508), .A2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n507), .A2(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G61), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n574), .A2(G86), .A3(new_n575), .A4(new_n520), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(G48), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n530), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n514), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n512), .A2(G92), .A3(new_n520), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n543), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n552), .A2(new_n599), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n595), .A2(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n467), .A2(new_n476), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT74), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n485), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n472), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n467), .A2(new_n472), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n614), .B(new_n622), .C1(G2100), .C2(new_n612), .ZN(G156));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT77), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n625), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT75), .B(KEYINPUT14), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n628), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(G401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT78), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n621), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1991), .B(G1996), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  MUX2_X1   g240(.A(new_n665), .B(new_n664), .S(new_n657), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT79), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n654), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n676), .A3(new_n654), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  NAND2_X1  g256(.A1(new_n485), .A2(G119), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n472), .A2(G107), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n684));
  INV_X1    g259(.A(G131), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n682), .B1(new_n683), .B2(new_n684), .C1(new_n685), .C2(new_n619), .ZN(new_n686));
  MUX2_X1   g261(.A(G25), .B(new_n686), .S(G29), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G24), .ZN(new_n690));
  INV_X1    g265(.A(G290), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT81), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT80), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n689), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n693), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT32), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1981), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT85), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1971), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT83), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n709), .B(new_n711), .Z(new_n712));
  AOI21_X1  g287(.A(new_n705), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n706), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n697), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n700), .B2(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT86), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(KEYINPUT86), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(KEYINPUT87), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n701), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n701), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT95), .B(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G26), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n489), .A2(G140), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n485), .A2(G128), .ZN(new_n735));
  OR2_X1    g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n736), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n731), .B1(new_n741), .B2(G34), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n480), .A2(new_n731), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  AOI22_X1  g320(.A1(G2067), .A2(new_n740), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n730), .B(new_n746), .C1(G2067), .C2(new_n740), .ZN(new_n747));
  NAND2_X1  g322(.A1(G164), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G27), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n758), .B1(new_n731), .B2(new_n620), .C1(new_n744), .C2(new_n745), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n747), .A2(new_n751), .A3(new_n752), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n476), .A2(G105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT92), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n763), .B(new_n765), .C1(G129), .C2(new_n485), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n489), .A2(G141), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT91), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n731), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G32), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n770), .A2(KEYINPUT94), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(KEYINPUT94), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n773), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n731), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G139), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n619), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G115), .A2(G2104), .ZN(new_n785));
  INV_X1    g360(.A(G127), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n488), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n472), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n777), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n775), .A2(new_n776), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n731), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n731), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  NOR2_X1   g377(.A1(G4), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n596), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n801), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n701), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT23), .ZN(new_n808));
  INV_X1    g383(.A(G299), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n701), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n804), .B2(G1348), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n760), .A2(new_n795), .A3(new_n806), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n799), .A2(new_n796), .A3(new_n800), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n815));
  NOR2_X1   g390(.A1(G5), .A2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G301), .B2(new_n701), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n814), .A2(new_n815), .B1(G1961), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n792), .A2(new_n793), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT90), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n701), .A2(G19), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n553), .B2(new_n701), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1341), .Z(new_n827));
  OAI221_X1 g402(.A(new_n827), .B1(G1961), .B2(new_n820), .C1(new_n814), .C2(new_n815), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n813), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n723), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n726), .A2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n723), .A2(new_n725), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n833), .B(new_n829), .C1(new_n723), .C2(new_n830), .ZN(G150));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n552), .A2(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n552), .A2(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n543), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT99), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n514), .B1(new_n841), .B2(KEYINPUT99), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n530), .A2(G93), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  INV_X1    g422(.A(new_n518), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n838), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n836), .A2(new_n850), .A3(new_n837), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n595), .A2(new_n603), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n857), .A3(new_n853), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n835), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n850), .A2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(G145));
  XOR2_X1   g448(.A(KEYINPUT104), .B(G37), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n739), .B(new_n505), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n791), .ZN(new_n877));
  INV_X1    g452(.A(new_n769), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n686), .B(new_n610), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n489), .A2(G142), .B1(G130), .B2(new_n485), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  INV_X1    g457(.A(G118), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n882), .A2(KEYINPUT102), .B1(new_n883), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(KEYINPUT102), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n880), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n480), .B(new_n620), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n879), .A2(new_n887), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n889), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n875), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n892), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n893), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n898), .A3(new_n888), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n900), .B(new_n897), .C1(new_n889), .C2(new_n888), .ZN(new_n906));
  INV_X1    g481(.A(new_n895), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n874), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n905), .A2(new_n910), .ZN(G395));
  XNOR2_X1  g486(.A(new_n606), .B(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n854), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n606), .B(KEYINPUT106), .Z(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n853), .A3(new_n852), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n596), .A2(new_n809), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n595), .A2(G299), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT41), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT108), .B1(new_n920), .B2(KEYINPUT41), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n920), .B(KEYINPUT107), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n913), .B2(new_n915), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G305), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G288), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(KEYINPUT109), .ZN(new_n934));
  MUX2_X1   g509(.A(new_n931), .B(new_n933), .S(new_n934), .Z(new_n935));
  INV_X1    g510(.A(new_n929), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n913), .B(new_n915), .C1(new_n924), .C2(new_n925), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n930), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n930), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n851), .A2(new_n599), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(G331));
  XNOR2_X1  g520(.A(G168), .B(G301), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n852), .A2(new_n853), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n852), .B2(new_n853), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n947), .A2(new_n948), .B1(new_n924), .B2(new_n925), .ZN(new_n949));
  INV_X1    g524(.A(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n854), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n920), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n852), .A2(new_n853), .A3(new_n946), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n935), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n949), .A2(new_n954), .A3(new_n935), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT43), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n921), .B(new_n923), .C1(new_n947), .C2(new_n948), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(new_n928), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n956), .ZN(new_n962));
  AND4_X1   g537(.A1(KEYINPUT43), .A2(new_n962), .A3(new_n958), .A4(new_n874), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n957), .B2(new_n958), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n966), .A2(new_n962), .A3(new_n958), .A4(new_n874), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(G397));
  INV_X1    g545(.A(KEYINPUT122), .ZN(new_n971));
  INV_X1    g546(.A(G1956), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n472), .B1(new_n468), .B2(new_n469), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT110), .B(G40), .Z(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n478), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n495), .B2(new_n504), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g553(.A(KEYINPUT50), .B(G1384), .C1(new_n495), .C2(new_n504), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n492), .A2(new_n494), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n498), .A2(new_n503), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n485), .A2(G126), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT56), .B(G2072), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n988), .A2(new_n975), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n809), .B2(KEYINPUT118), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n994));
  NAND3_X1  g569(.A1(G299), .A2(new_n994), .A3(KEYINPUT57), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n980), .A2(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT61), .B1(new_n996), .B2(KEYINPUT120), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n995), .ZN(new_n998));
  INV_X1    g573(.A(new_n974), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n471), .A2(new_n479), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n976), .A2(new_n977), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1956), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n975), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n987), .B(G1384), .C1(new_n495), .C2(new_n504), .ZN(new_n1005));
  INV_X1    g580(.A(new_n990), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n998), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n980), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n997), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n802), .B1(new_n978), .B2(new_n979), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n976), .A2(new_n975), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(G2067), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1014), .A2(new_n1016), .A3(new_n595), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n595), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT60), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1004), .A2(G1996), .A3(new_n1005), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT58), .B(G1341), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n553), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1015), .A2(G2067), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n975), .A3(new_n1002), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1028), .B2(new_n802), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1024), .A2(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n1010), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1033));
  OAI211_X1 g608(.A(new_n553), .B(new_n1033), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1019), .A2(new_n1031), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1012), .B1(new_n997), .B2(new_n1011), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1013), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1010), .B1(new_n996), .B2(new_n1018), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n971), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n975), .C1(new_n976), .C2(KEYINPUT45), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1043), .A3(new_n989), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n729), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT115), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1027), .A2(new_n745), .A3(new_n975), .A4(new_n1002), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1001), .A2(KEYINPUT116), .A3(new_n745), .A4(new_n1002), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(new_n1052), .A3(new_n729), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1046), .A2(new_n1051), .A3(G168), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(KEYINPUT123), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  INV_X1    g633(.A(new_n729), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1005), .B1(new_n1004), .B2(KEYINPUT114), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1043), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1061), .A2(new_n1052), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1055), .B1(new_n1062), .B2(new_n1046), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G286), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1065), .A3(new_n1056), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1027), .A2(new_n796), .A3(new_n975), .A4(new_n1002), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n978), .A2(G2090), .A3(new_n979), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1070), .B(G8), .C1(new_n1072), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n579), .A2(new_n582), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n514), .B1(new_n576), .B2(new_n577), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n580), .A2(new_n581), .ZN(new_n1082));
  OAI21_X1  g657(.A(G1981), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1015), .A2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1055), .B1(new_n976), .B2(new_n975), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n708), .A2(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1091), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1068), .B(KEYINPUT55), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1074), .A2(new_n1071), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1055), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1078), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n988), .A2(new_n750), .A3(new_n975), .A4(new_n989), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1028), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(G2078), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(G40), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n988), .A2(G160), .A3(new_n989), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1108), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT124), .B1(new_n1114), .B2(G171), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1060), .A2(new_n1043), .A3(new_n1111), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1107), .A2(new_n1106), .B1(new_n1028), .B2(new_n1109), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(G301), .A4(new_n1113), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1078), .A2(new_n1100), .A3(new_n1125), .A4(new_n1103), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1114), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1119), .A2(KEYINPUT126), .A3(new_n1113), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(G171), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(G301), .A3(new_n1116), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(KEYINPUT54), .A3(new_n1131), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1105), .A2(new_n1124), .A3(new_n1126), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n997), .A2(new_n1011), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1019), .A2(new_n1032), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n997), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(KEYINPUT122), .A3(new_n1038), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1040), .A2(new_n1067), .A3(new_n1133), .A4(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1091), .A2(new_n1097), .A3(new_n708), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1080), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1093), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1091), .A2(new_n1099), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1078), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n988), .A2(new_n975), .A3(new_n989), .ZN(new_n1148));
  AOI22_X1  g723(.A1(KEYINPUT112), .A2(new_n1071), .B1(new_n1148), .B2(new_n1073), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1055), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1145), .B1(new_n1151), .B2(new_n1070), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  OAI21_X1  g728(.A(G8), .B1(new_n1077), .B2(new_n1072), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1101), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1152), .A2(new_n1155), .A3(new_n1063), .A4(G168), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1152), .A2(new_n1063), .A3(G168), .A4(new_n1103), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1147), .A2(new_n1156), .B1(new_n1157), .B2(new_n1153), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1156), .A2(new_n1147), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1146), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1161));
  AND4_X1   g736(.A1(G171), .A2(new_n1105), .A3(new_n1117), .A4(new_n1126), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1058), .A2(new_n1163), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1141), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n988), .A2(new_n1000), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1168), .A2(G1986), .A3(G290), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n691), .A2(new_n673), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT111), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n738), .B(G2067), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n878), .A2(G1996), .ZN(new_n1174));
  INV_X1    g749(.A(G1996), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n769), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n686), .B(new_n688), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1168), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1166), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1182));
  AND2_X1   g757(.A1(new_n1169), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1169), .A2(new_n1182), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1167), .B1(new_n769), .B2(new_n1173), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1168), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT46), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1167), .B2(new_n1175), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1186), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  INV_X1    g766(.A(new_n688), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n686), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1177), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n738), .A2(G2067), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1185), .B(new_n1191), .C1(new_n1167), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1181), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g773(.A1(new_n967), .A2(new_n968), .ZN(new_n1200));
  NOR3_X1   g774(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n680), .B(new_n1201), .C1(new_n908), .C2(new_n903), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1202), .ZN(G308));
  NAND2_X1  g777(.A1(new_n896), .A2(new_n904), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n680), .A2(new_n1201), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n1204), .B(new_n1205), .C1(new_n967), .C2(new_n968), .ZN(G225));
endmodule


