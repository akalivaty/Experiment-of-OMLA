//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n202), .A2(G77), .A3(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n204), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n227), .A2(G1), .A3(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n205), .A2(G50), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n211), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT0), .Z(new_n236));
  NOR4_X1   g0036(.A1(new_n223), .A2(new_n224), .A3(new_n233), .A4(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT75), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT10), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n255), .A2(KEYINPUT10), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n260), .B1(new_n261), .B2(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n226), .B2(new_n228), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT70), .B1(new_n265), .B2(new_n225), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n268), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT69), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n269), .B2(new_n273), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n274), .A2(new_n277), .B1(new_n279), .B2(G226), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n267), .A2(G190), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT74), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  AND4_X1   g0085(.A1(new_n226), .A2(new_n228), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G50), .B1(new_n231), .B2(G1), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G50), .ZN(new_n289));
  INV_X1    g0089(.A(new_n284), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n231), .A2(new_n292), .A3(KEYINPUT71), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G20), .B2(G33), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n203), .A2(KEYINPUT8), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT8), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G58), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n231), .A2(G33), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n296), .A2(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n205), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n231), .B1(new_n201), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n226), .A2(new_n228), .A3(new_n285), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n291), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT9), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n267), .A2(new_n280), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT9), .B(new_n291), .C1(new_n307), .C2(new_n308), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n256), .B(new_n257), .C1(new_n283), .C2(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n281), .B(KEYINPUT74), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n255), .A4(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(new_n309), .C1(G179), .C2(new_n312), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT72), .B(G107), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n258), .B2(new_n326), .C1(new_n262), .C2(new_n213), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n266), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n277), .A2(new_n274), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  INV_X1    g0130(.A(new_n279), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n320), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n331), .B2(new_n330), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n266), .B2(new_n327), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n226), .A2(new_n228), .A3(new_n285), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n231), .A2(G1), .ZN(new_n339));
  NOR4_X1   g0139(.A1(new_n338), .A2(new_n290), .A3(new_n261), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G20), .A2(G77), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n303), .B2(new_n343), .C1(new_n296), .C2(new_n302), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n338), .B1(new_n261), .B2(new_n290), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n333), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n335), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n341), .B(new_n345), .C1(new_n332), .C2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n324), .B(new_n347), .C1(new_n349), .C2(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n225), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n354));
  OAI211_X1 g0154(.A(G232), .B(new_n276), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT79), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n279), .A2(new_n357), .A3(G232), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G33), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n362), .A3(G223), .A4(new_n259), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n360), .A2(new_n362), .A3(G226), .A4(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n266), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n266), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n359), .A2(new_n329), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT80), .B1(new_n371), .B2(G179), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n258), .A2(new_n373), .A3(G20), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n360), .A2(new_n362), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n375), .B2(new_n231), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n293), .B2(new_n295), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n231), .B1(new_n205), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT77), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n205), .A2(new_n380), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G20), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT77), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n296), .C2(new_n378), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n382), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n373), .B1(new_n258), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n204), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n293), .A2(new_n295), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G159), .B1(new_n383), .B2(G20), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n388), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n395), .A3(new_n338), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n302), .A2(new_n339), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n286), .B1(new_n290), .B2(new_n302), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n357), .B1(new_n279), .B2(G232), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n329), .B(new_n367), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n320), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n366), .A2(new_n266), .A3(new_n369), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n369), .B1(new_n366), .B2(new_n266), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n356), .A2(new_n358), .B1(new_n274), .B2(new_n277), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT80), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n336), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n372), .A2(new_n399), .A3(new_n403), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n409), .A2(new_n403), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n399), .A4(new_n372), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n396), .A2(new_n398), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n407), .A3(new_n350), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n402), .A2(new_n348), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT17), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n414), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n296), .A2(new_n289), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n303), .A2(new_n261), .B1(new_n231), .B2(G68), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n338), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT11), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n339), .A2(new_n204), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n284), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT12), .B1(new_n284), .B2(G68), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n286), .A2(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n274), .A2(new_n277), .B1(new_n279), .B2(G238), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n360), .A2(new_n362), .A3(G232), .A4(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n360), .A2(new_n362), .A3(G226), .A4(new_n259), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G97), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n266), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n436), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n279), .A2(G238), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n329), .A2(new_n442), .A3(new_n436), .A4(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n446), .B2(G169), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n435), .B(G169), .C1(new_n443), .C2(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n437), .A2(new_n442), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT13), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(new_n436), .A3(new_n442), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(G179), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n434), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(G200), .ZN(new_n455));
  INV_X1    g0255(.A(new_n434), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(G190), .A3(new_n451), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n352), .A2(new_n423), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n258), .A2(G257), .A3(new_n259), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n375), .A2(G303), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n266), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n269), .A2(new_n273), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(G274), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n269), .A2(new_n273), .B1(new_n469), .B2(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G270), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n275), .A2(G33), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n286), .A2(G116), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n290), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(G33), .B2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n292), .A2(G97), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(G20), .B2(new_n476), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(new_n338), .A3(KEYINPUT20), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n480), .B2(new_n338), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n473), .A2(new_n483), .A3(KEYINPUT21), .A4(G169), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n472), .A2(new_n470), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(new_n483), .A3(G179), .A4(new_n465), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n473), .A2(new_n483), .A3(G169), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n483), .B1(new_n473), .B2(G200), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n350), .B2(new_n473), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n468), .A2(new_n215), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n353), .B2(new_n354), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n292), .A2(new_n476), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G238), .A2(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n330), .B2(G1698), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n258), .ZN(new_n499));
  INV_X1    g0299(.A(new_n266), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n466), .A2(G274), .A3(new_n468), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n330), .A2(G1698), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G238), .B2(G1698), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n505), .A2(new_n375), .B1(new_n292), .B2(new_n476), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n266), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n274), .A2(new_n468), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(G179), .A4(new_n495), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n360), .A2(new_n362), .A3(new_n231), .A4(G68), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n303), .A2(new_n207), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(KEYINPUT19), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(G87), .A2(G97), .ZN(new_n514));
  NAND3_X1  g0314(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n326), .A2(new_n514), .B1(new_n231), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n338), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT15), .B(G87), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n343), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n286), .A2(new_n519), .A3(new_n474), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n343), .A2(new_n290), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n517), .A2(new_n522), .A3(KEYINPUT84), .A4(new_n523), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n510), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n517), .A2(new_n523), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n286), .A2(new_n474), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G87), .ZN(new_n533));
  OAI21_X1  g0333(.A(G200), .B1(new_n501), .B2(new_n502), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n507), .A2(new_n508), .A3(G190), .A4(new_n495), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n530), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT85), .B1(new_n528), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n360), .A2(new_n362), .A3(G244), .A4(new_n259), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G283), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n266), .B1(G257), .B2(new_n471), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n470), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n320), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n336), .A3(new_n470), .ZN(new_n550));
  XOR2_X1   g0350(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n551));
  NAND2_X1  g0351(.A1(new_n208), .A2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n209), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(G20), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n392), .A2(G77), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n326), .B1(new_n389), .B2(new_n390), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n338), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n290), .A2(KEYINPUT82), .A3(new_n207), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n284), .B2(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n531), .B2(new_n207), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n549), .A2(new_n550), .A3(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n561), .A2(new_n567), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n548), .A2(G200), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n547), .A2(G190), .A3(new_n470), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n360), .A2(new_n362), .A3(G257), .A4(G1698), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n360), .A2(new_n362), .A3(G250), .A4(new_n259), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n266), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n469), .A2(new_n468), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n466), .A2(G264), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n470), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n578), .A2(new_n470), .A3(G179), .A4(new_n580), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n208), .A2(G20), .ZN(new_n585));
  OAI22_X1  g0385(.A1(KEYINPUT23), .A2(new_n585), .B1(new_n303), .B2(new_n476), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n326), .A2(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT23), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n360), .A2(new_n362), .A3(new_n231), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n258), .A2(new_n591), .A3(new_n231), .A4(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n588), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n308), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G13), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G1), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(G20), .A3(new_n208), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT25), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n532), .A2(G107), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n584), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n578), .A2(new_n470), .A3(new_n350), .A4(new_n580), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n578), .A2(new_n470), .A3(new_n580), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n597), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n596), .B1(new_n588), .B2(new_n593), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n338), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n613), .A3(new_n605), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n569), .A2(new_n573), .A3(new_n607), .A4(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n460), .A2(new_n493), .A3(new_n539), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT86), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n510), .A2(new_n524), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n548), .A2(new_n320), .B1(new_n561), .B2(new_n567), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(new_n536), .A3(new_n550), .A4(new_n618), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n528), .A2(new_n536), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n536), .ZN(new_n625));
  INV_X1    g0425(.A(new_n569), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n621), .B1(KEYINPUT26), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n490), .A2(new_n486), .A3(new_n484), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n613), .A2(new_n605), .B1(new_n582), .B2(new_n583), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n629), .A2(KEYINPUT87), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n534), .A2(new_n535), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n529), .B1(G87), .B2(new_n532), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n633), .B1(new_n510), .B2(new_n524), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n573), .A2(new_n634), .A3(new_n569), .A4(new_n614), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n487), .A2(new_n490), .A3(new_n607), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n631), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n628), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n460), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n421), .A2(new_n422), .ZN(new_n642));
  INV_X1    g0442(.A(new_n347), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n458), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n454), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n411), .A2(new_n414), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n316), .B(new_n319), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n322), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n600), .A2(new_n231), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n483), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n493), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n487), .B2(new_n490), .ZN(new_n658));
  OAI21_X1  g0458(.A(G330), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n655), .B1(new_n598), .B2(new_n606), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n607), .A2(new_n660), .A3(new_n614), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n607), .A2(new_n660), .A3(new_n614), .A4(KEYINPUT88), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  INV_X1    g0465(.A(new_n655), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n607), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n630), .A2(KEYINPUT89), .A3(new_n655), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n663), .A2(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n630), .A2(new_n666), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n655), .B1(new_n487), .B2(new_n490), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n670), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n234), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n326), .A2(new_n476), .A3(new_n514), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n232), .B2(new_n678), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n620), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n537), .A2(new_n538), .A3(new_n569), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  INV_X1    g0488(.A(new_n618), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n636), .B2(new_n637), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT90), .B1(new_n691), .B2(new_n666), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n685), .B1(new_n627), .B2(new_n684), .ZN(new_n693));
  INV_X1    g0493(.A(new_n637), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n618), .B1(new_n694), .B2(new_n635), .ZN(new_n695));
  OAI211_X1 g0495(.A(KEYINPUT90), .B(new_n666), .C1(new_n693), .C2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT29), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n655), .B1(new_n628), .B2(new_n639), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n501), .A2(new_n502), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n547), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n473), .A2(new_n336), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n609), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n609), .A2(new_n547), .A3(new_n704), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n485), .A2(G179), .A3(new_n465), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n704), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n548), .A3(new_n473), .A4(new_n581), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n714), .B2(new_n655), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n615), .A2(new_n539), .A3(new_n493), .A4(new_n666), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n703), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n702), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n683), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n599), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n275), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n677), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n230), .B1(G20), .B2(new_n320), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n676), .A2(new_n375), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G355), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G116), .B2(new_n234), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n250), .A2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n232), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n258), .B(new_n676), .C1(new_n738), .C2(new_n467), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n727), .B1(new_n733), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n231), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n350), .A3(G200), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n258), .B1(new_n743), .B2(new_n208), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n231), .A2(new_n336), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n231), .A2(new_n336), .A3(KEYINPUT92), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n350), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n744), .B1(new_n753), .B2(G58), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n742), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n378), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n750), .A2(new_n755), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n754), .B(new_n758), .C1(new_n261), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n745), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n204), .B1(new_n764), .B2(new_n214), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n751), .A2(new_n336), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n207), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n761), .A2(new_n350), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n289), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n760), .A2(new_n765), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT93), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n753), .A2(G322), .B1(new_n762), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  INV_X1    g0577(.A(new_n764), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n770), .A2(G326), .B1(new_n778), .B2(G303), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n743), .ZN(new_n781));
  INV_X1    g0581(.A(new_n756), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n258), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n783), .B1(new_n784), .B2(new_n768), .C1(new_n759), .C2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n777), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n774), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT95), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n728), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n741), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n657), .A2(new_n658), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n731), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n703), .ZN(new_n798));
  INV_X1    g0598(.A(new_n727), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n798), .A2(new_n659), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n346), .A2(new_n655), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n351), .B2(new_n349), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n347), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n643), .A2(new_n666), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n699), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n699), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n727), .B1(new_n812), .B2(new_n720), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n720), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n728), .A2(new_n729), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n799), .B1(new_n815), .B2(new_n261), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n258), .B(new_n769), .C1(G311), .C2(new_n782), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n476), .B2(new_n759), .C1(new_n784), .C2(new_n752), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n214), .A2(new_n743), .B1(new_n764), .B2(new_n208), .ZN(new_n819));
  INV_X1    g0619(.A(G303), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n763), .A2(new_n780), .B1(new_n771), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n762), .A2(G150), .B1(new_n770), .B2(G137), .ZN(new_n823));
  INV_X1    g0623(.A(G143), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n752), .B2(new_n824), .C1(new_n378), .C2(new_n759), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n258), .B1(new_n756), .B2(new_n829), .C1(new_n768), .C2(new_n203), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT97), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n289), .A2(new_n764), .B1(new_n743), .B2(new_n204), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n822), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n816), .B1(new_n836), .B2(new_n791), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT98), .Z(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n730), .B2(new_n809), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n814), .A2(new_n839), .ZN(G384));
  NOR2_X1   g0640(.A1(new_n724), .A2(new_n275), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  INV_X1    g0642(.A(new_n653), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n399), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n423), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n410), .A2(new_n419), .A3(new_n844), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n410), .A2(new_n419), .A3(new_n849), .A4(new_n844), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n850), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n387), .A2(new_n338), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n389), .A2(new_n390), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G68), .B1(new_n393), .B2(new_n385), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n858), .B2(new_n382), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n398), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n415), .A2(new_n418), .B1(new_n860), .B2(new_n843), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(new_n372), .A3(new_n403), .A4(new_n409), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT100), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n843), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(new_n419), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n850), .ZN(new_n869));
  INV_X1    g0669(.A(new_n865), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n423), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n864), .A2(new_n869), .A3(new_n871), .A4(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n854), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n434), .A2(new_n655), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT99), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n454), .A2(new_n458), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n454), .A2(new_n458), .A3(KEYINPUT99), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n447), .A2(new_n453), .A3(new_n874), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n874), .A2(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n714), .A2(new_n655), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT31), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n881), .A4(new_n655), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n718), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n879), .A2(new_n886), .A3(new_n809), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n842), .B1(new_n873), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n879), .A2(new_n886), .A3(new_n842), .A4(new_n809), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n864), .A2(new_n869), .A3(new_n871), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n853), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n872), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT103), .Z(new_n894));
  AND2_X1   g0694(.A1(new_n460), .A2(new_n886), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n703), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(new_n807), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n699), .B2(new_n809), .ZN(new_n899));
  INV_X1    g0699(.A(new_n879), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n872), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n646), .B2(new_n653), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n891), .B2(new_n872), .ZN(new_n905));
  XOR2_X1   g0705(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n906));
  AND3_X1   g0706(.A1(new_n854), .A2(new_n872), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n454), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n666), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n903), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n698), .A2(new_n460), .A3(new_n701), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(new_n648), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n911), .B(new_n913), .Z(new_n914));
  AOI21_X1  g0714(.A(new_n841), .B1(new_n897), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n897), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n230), .A2(new_n231), .A3(new_n476), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n553), .A2(new_n556), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT36), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n738), .A2(G77), .A3(new_n380), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n204), .B2(new_n202), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n599), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n916), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI22_X1  g0726(.A1(new_n763), .A2(new_n378), .B1(new_n771), .B2(new_n824), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n768), .A2(new_n204), .B1(new_n764), .B2(new_n203), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n759), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n202), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n753), .A2(G150), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n743), .A2(new_n261), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n375), .B(new_n933), .C1(G137), .C2(new_n782), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n929), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n759), .A2(new_n780), .B1(new_n326), .B2(new_n768), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT111), .Z(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n375), .B1(new_n756), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n771), .A2(new_n785), .B1(new_n743), .B2(new_n207), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(G294), .C2(new_n762), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT46), .B1(new_n778), .B2(G116), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n753), .B2(G303), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n935), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n728), .ZN(new_n948));
  INV_X1    g0748(.A(new_n732), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n676), .B2(new_n518), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n676), .A2(new_n258), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n246), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n799), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n634), .B1(new_n633), .B2(new_n666), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n618), .A2(new_n633), .A3(new_n666), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n948), .B(new_n953), .C1(new_n796), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n663), .A2(new_n664), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n667), .A2(new_n668), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n672), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n493), .A2(new_n656), .ZN(new_n962));
  INV_X1    g0762(.A(new_n658), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n703), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n669), .A2(new_n673), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI221_X4 g0766(.A(new_n672), .B1(new_n667), .B2(new_n668), .C1(new_n663), .C2(new_n664), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n673), .B1(new_n958), .B2(new_n959), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n659), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT29), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n666), .B1(new_n693), .B2(new_n695), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT90), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n971), .B1(new_n974), .B2(new_n696), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n970), .B(new_n720), .C1(new_n975), .C2(new_n700), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT108), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n573), .B(new_n569), .C1(new_n570), .C2(new_n666), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n626), .A2(new_n655), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n674), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n674), .A2(new_n983), .A3(KEYINPUT44), .A4(new_n981), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n979), .A2(new_n980), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n671), .A4(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n671), .B(new_n990), .C1(new_n669), .C2(new_n673), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n991), .A2(new_n994), .B1(KEYINPUT109), .B2(new_n670), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n989), .B1(new_n988), .B2(new_n995), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n721), .B1(new_n978), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n677), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(new_n725), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT105), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n981), .A2(KEYINPUT104), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT104), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n990), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n607), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1002), .B1(new_n1006), .B2(new_n626), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n990), .B(KEYINPUT104), .ZN(new_n1008));
  OAI211_X1 g0808(.A(KEYINPUT105), .B(new_n569), .C1(new_n1008), .C2(new_n607), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1009), .A3(new_n666), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n968), .A2(new_n990), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n956), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1008), .A2(new_n659), .A3(new_n669), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1010), .A2(new_n1016), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT110), .B1(new_n1001), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n976), .A2(KEYINPUT108), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n702), .A2(new_n977), .A3(new_n720), .A4(new_n970), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n997), .C2(new_n996), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1000), .B1(new_n1028), .B2(new_n722), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1024), .B(KEYINPUT110), .C1(new_n1029), .C2(new_n726), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n957), .B1(new_n1025), .B2(new_n1031), .ZN(G387));
  NAND2_X1  g0832(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n677), .C1(new_n722), .C2(new_n970), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n734), .A2(new_n679), .B1(new_n208), .B2(new_n676), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n243), .A2(new_n467), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n680), .B(new_n467), .C1(new_n204), .C2(new_n261), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n301), .A2(new_n289), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n951), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n733), .B1(new_n1041), .B2(KEYINPUT112), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT112), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n727), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n519), .A2(new_n521), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n767), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n289), .B2(new_n752), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT113), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n778), .A2(G77), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G159), .A2(new_n770), .B1(new_n762), .B2(new_n301), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n258), .B1(new_n756), .B2(new_n297), .C1(new_n207), .C2(new_n743), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n930), .B2(G68), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n258), .B1(new_n782), .B2(G326), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n768), .A2(new_n780), .B1(new_n764), .B2(new_n784), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n762), .A2(G311), .B1(new_n770), .B2(G322), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n752), .B2(new_n938), .C1(new_n820), .C2(new_n759), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1054), .B1(new_n476), .B2(new_n743), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1053), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT114), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n791), .B1(new_n1064), .B2(KEYINPUT114), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1044), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n669), .A2(new_n731), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(new_n1068), .B1(new_n726), .B2(new_n970), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1034), .A2(new_n1069), .ZN(G393));
  AOI21_X1  g0870(.A(new_n949), .B1(G97), .B2(new_n676), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n253), .A2(new_n951), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n799), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n258), .B1(new_n756), .B2(new_n824), .C1(new_n214), .C2(new_n743), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n768), .A2(new_n261), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n202), .B2(new_n762), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n204), .B2(new_n764), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1074), .B(new_n1077), .C1(new_n301), .C2(new_n930), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n752), .A2(new_n378), .B1(new_n297), .B2(new_n771), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n763), .A2(new_n820), .B1(new_n768), .B2(new_n476), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n258), .B1(new_n782), .B2(G322), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n208), .B2(new_n743), .C1(new_n759), .C2(new_n784), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G283), .C2(new_n778), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n752), .A2(new_n785), .B1(new_n938), .B2(new_n771), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1078), .A2(new_n1080), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1073), .B1(new_n1087), .B2(new_n791), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1008), .B2(new_n731), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n998), .B2(new_n726), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n978), .A2(new_n998), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1028), .A2(new_n677), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(G390));
  OAI21_X1  g0893(.A(new_n910), .B1(new_n899), .B2(new_n900), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n974), .A2(new_n696), .A3(new_n807), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n806), .A3(new_n879), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n873), .A2(new_n910), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n908), .A2(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n703), .B1(new_n885), .B2(new_n718), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n879), .A3(new_n809), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT115), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n854), .A2(new_n872), .A3(new_n906), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1094), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1096), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT115), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1100), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n719), .A2(new_n809), .A3(new_n879), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1098), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1101), .A2(new_n726), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n908), .A2(new_n729), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n799), .B1(new_n815), .B2(new_n302), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n375), .B1(new_n756), .B2(new_n784), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G87), .B2(new_n778), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n752), .B2(new_n476), .C1(new_n207), .C2(new_n759), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n743), .A2(new_n204), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n780), .A2(new_n771), .B1(new_n763), .B2(new_n326), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1075), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n753), .A2(G132), .B1(G128), .B2(new_n770), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n258), .B1(new_n756), .B2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n768), .A2(new_n378), .B1(new_n201), .B2(new_n743), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G137), .C2(new_n762), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n778), .A2(G150), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT53), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI22_X1  g0932(.A1(new_n930), .A2(new_n1132), .B1(KEYINPUT53), .B2(new_n1130), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1125), .A2(new_n1129), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1123), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1114), .B(new_n1115), .C1(new_n791), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1113), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1101), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n460), .A2(new_n1099), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n912), .A2(new_n648), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n879), .B1(new_n1099), .B2(new_n809), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1110), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1095), .A2(new_n806), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n899), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n703), .B(new_n808), .C1(new_n717), .C2(new_n718), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1100), .B1(new_n1146), .B2(new_n879), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1143), .A2(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n678), .B1(new_n1139), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1101), .A2(new_n1112), .A3(new_n1109), .A4(new_n1149), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1138), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1141), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(G330), .B1(new_n888), .B2(new_n892), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n323), .A2(new_n309), .A3(new_n843), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n309), .A2(new_n843), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n316), .A2(new_n319), .A3(new_n322), .A4(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1161), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT119), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1158), .A3(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1157), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(G330), .C1(new_n888), .C2(new_n892), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1173), .A2(new_n911), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n911), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1156), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n911), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n911), .A2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1174), .A3(new_n1173), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1152), .A2(new_n1155), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1179), .B(new_n677), .C1(KEYINPUT57), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n725), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n930), .A2(new_n1045), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n207), .B2(new_n763), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT118), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n258), .A2(G41), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n780), .B2(new_n756), .C1(new_n768), .C2(new_n204), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1049), .B1(new_n203), .B2(new_n743), .C1(new_n771), .C2(new_n476), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G107), .C2(new_n753), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1191), .A2(KEYINPUT58), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n930), .A2(G137), .B1(new_n753), .B2(G128), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n770), .A2(G125), .B1(new_n767), .B2(G150), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n762), .A2(G132), .B1(new_n778), .B2(new_n1132), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  INV_X1    g1003(.A(G41), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n292), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n782), .B2(G124), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n378), .B2(new_n743), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1202), .A2(new_n1203), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT58), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G50), .B(new_n1192), .C1(new_n292), .C2(new_n1204), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1197), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n791), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n815), .A2(new_n201), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n727), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(new_n1172), .C2(new_n729), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1187), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1186), .A2(new_n1217), .ZN(G375));
  NOR2_X1   g1018(.A1(new_n768), .A2(new_n289), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n771), .A2(new_n829), .B1(new_n764), .B2(new_n378), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n762), .C2(new_n1132), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n375), .B1(new_n782), .B2(G128), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n203), .B2(new_n743), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n753), .B2(G137), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1221), .B(new_n1224), .C1(new_n297), .C2(new_n759), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n326), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n930), .A2(new_n1226), .B1(new_n753), .B2(G283), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n763), .A2(new_n476), .B1(new_n764), .B2(new_n207), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G294), .B2(new_n770), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n258), .B(new_n933), .C1(G303), .C2(new_n782), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1046), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1225), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n728), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n799), .B1(new_n815), .B2(new_n204), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n879), .C2(new_n730), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1148), .B2(new_n725), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1149), .A2(new_n1000), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G381));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1034), .A2(new_n802), .A3(new_n1241), .A4(new_n1069), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1244), .A2(new_n1245), .A3(G390), .A4(G381), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n957), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT110), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1028), .A2(new_n722), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1000), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n726), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1247), .B1(new_n1253), .B2(new_n1030), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1246), .A2(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(KEYINPUT122), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT122), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G375), .A2(G378), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(G407));
  INV_X1    g1059(.A(new_n1258), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G343), .C2(new_n1260), .ZN(G409));
  AOI21_X1  g1061(.A(new_n1153), .B1(new_n1186), .B2(new_n1217), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n654), .A2(G213), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1139), .A2(new_n1150), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n677), .A3(new_n1152), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1138), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1215), .B1(new_n1267), .B2(new_n726), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1185), .A2(new_n1250), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1262), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1236), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(new_n1238), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n677), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1241), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1276), .A2(new_n677), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1238), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1236), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT124), .B1(new_n1283), .B2(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G384), .B(new_n1273), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT123), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT123), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1288), .A3(G384), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NOR4_X1   g1094(.A1(new_n1262), .A2(new_n1271), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G387), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n957), .B(G390), .C1(new_n1025), .C2(new_n1031), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT126), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT127), .B1(new_n1254), .B2(G390), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1254), .A2(new_n1303), .A3(G390), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1299), .A2(new_n1301), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G396), .B(G393), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1254), .B2(G390), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1300), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G375), .A2(G378), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1185), .A2(new_n1250), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1315), .A2(new_n1316), .B1(G213), .B2(new_n654), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1263), .A2(KEYINPUT125), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1285), .A2(new_n1290), .A3(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1314), .A2(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1285), .A2(new_n1290), .A3(new_n1318), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1320), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1296), .A2(new_n1313), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1153), .A2(new_n1316), .A3(new_n1268), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1156), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1177), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n678), .B1(new_n1156), .B2(new_n1178), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1216), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1263), .B(new_n1327), .C1(new_n1332), .C2(new_n1153), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT62), .B1(new_n1333), .B2(new_n1291), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1285), .A2(new_n1290), .A3(new_n1320), .A4(new_n1318), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1324), .B(new_n1336), .C1(new_n1262), .C2(new_n1271), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1314), .A2(new_n1317), .A3(new_n1338), .A4(new_n1292), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1334), .A2(new_n1335), .A3(new_n1337), .A4(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1311), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1326), .A2(new_n1342), .ZN(G405));
  NAND3_X1  g1143(.A1(new_n1260), .A2(new_n1291), .A3(new_n1314), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1292), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1313), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1341), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


