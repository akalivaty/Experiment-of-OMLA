//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  XOR2_X1   g000(.A(G110), .B(G122), .Z(new_n187));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT3), .A2(G107), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT77), .A2(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT77), .A2(G104), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT3), .A2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n188), .B(G101), .C1(new_n192), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT3), .A2(G107), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(G104), .B2(new_n189), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n193), .A2(new_n194), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT77), .A2(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT77), .A2(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n207), .A2(KEYINPUT78), .A3(new_n188), .A4(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT2), .B(G113), .Z(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT67), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT67), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(G116), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n210), .B1(new_n217), .B2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(new_n210), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n207), .A2(G101), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n202), .A2(new_n206), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n209), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT5), .A3(new_n212), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT5), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(G113), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n217), .A2(new_n210), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n194), .B1(new_n204), .B2(new_n205), .ZN(new_n236));
  NAND2_X1  g050(.A1(G104), .A2(G107), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(G101), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT80), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n236), .A2(new_n240), .A3(G101), .A4(new_n237), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n226), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n228), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n209), .A2(new_n223), .A3(new_n227), .ZN(new_n245));
  INV_X1    g059(.A(new_n187), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n245), .B(new_n246), .C1(new_n235), .C2(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT0), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT0), .B(G128), .Z(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT75), .B(G125), .Z(new_n255));
  OR2_X1    g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT65), .B(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n249), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n258), .A2(new_n263), .A3(new_n264), .A4(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n255), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G224), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n187), .C1(new_n228), .C2(new_n243), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n248), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n248), .A2(new_n274), .A3(KEYINPUT84), .A4(new_n272), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n268), .B(KEYINPUT86), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n256), .ZN(new_n282));
  INV_X1    g096(.A(new_n271), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n271), .B2(KEYINPUT87), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n269), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n282), .A2(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n187), .B(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n239), .A2(new_n226), .A3(new_n241), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n234), .B2(new_n233), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n243), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n247), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n279), .A2(new_n280), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n277), .B2(new_n278), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n297), .A3(new_n295), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n301), .A2(KEYINPUT88), .A3(new_n297), .A4(new_n295), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT89), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n303), .A2(new_n304), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n198), .A2(new_n199), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n225), .B1(new_n202), .B2(new_n206), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT78), .B1(new_n313), .B2(new_n188), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n254), .B(new_n227), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n209), .A2(KEYINPUT79), .A3(new_n254), .A4(new_n227), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G134), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G137), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(G137), .ZN(new_n323));
  INV_X1    g137(.A(G137), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT11), .A3(G134), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT64), .A2(G131), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n322), .A2(new_n325), .A3(new_n327), .A4(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(KEYINPUT68), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n251), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n265), .B1(new_n337), .B2(new_n249), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n239), .A2(new_n226), .A3(new_n241), .A4(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(KEYINPUT81), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(KEYINPUT81), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n242), .A2(new_n336), .A3(new_n267), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n319), .A2(new_n335), .A3(new_n342), .A4(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n242), .A2(new_n267), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n292), .A2(new_n347), .A3(new_n338), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(KEYINPUT81), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n351));
  INV_X1    g165(.A(new_n331), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n242), .A2(new_n267), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n340), .B2(new_n341), .ZN(new_n355));
  INV_X1    g169(.A(new_n335), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT12), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n345), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  INV_X1    g173(.A(G227), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G953), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n359), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n342), .A2(new_n344), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n313), .A2(new_n188), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n200), .A2(new_n208), .B1(new_n366), .B2(new_n226), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT79), .B1(new_n367), .B2(new_n254), .ZN(new_n368));
  INV_X1    g182(.A(new_n318), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT82), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n348), .A2(new_n349), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n343), .B1(new_n372), .B2(new_n336), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n319), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n335), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n345), .A2(new_n362), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n364), .B(G469), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(G469), .A2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n345), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n363), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n377), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n351), .B1(new_n350), .B2(new_n335), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n355), .A2(KEYINPUT12), .A3(new_n331), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n380), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT9), .B(G234), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G221), .B1(new_n392), .B2(G902), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n311), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  AOI211_X1 g209(.A(G469), .B(G902), .C1(new_n382), .C2(new_n387), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT83), .B(new_n393), .C1(new_n396), .C2(new_n380), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n308), .A2(new_n310), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  INV_X1    g215(.A(G953), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G210), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n400), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT26), .B(G101), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n333), .A2(new_n254), .A3(new_n334), .ZN(new_n407));
  INV_X1    g221(.A(new_n223), .ZN(new_n408));
  INV_X1    g222(.A(new_n323), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n321), .A2(G137), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G131), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n322), .A2(new_n325), .A3(new_n412), .A4(new_n323), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n411), .B(new_n413), .C1(new_n261), .C2(new_n266), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT28), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n331), .A2(new_n254), .ZN(new_n417));
  INV_X1    g231(.A(new_n414), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n223), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n406), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n417), .B2(new_n418), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n423), .A3(new_n223), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(KEYINPUT70), .A3(new_n415), .A4(new_n406), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT31), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G472), .A2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n399), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n416), .A2(new_n419), .ZN(new_n433));
  INV_X1    g247(.A(new_n406), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n425), .A2(new_n426), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT32), .A3(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n430), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n432), .A2(new_n439), .B1(new_n440), .B2(KEYINPUT71), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n440), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n442));
  INV_X1    g256(.A(G472), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n407), .A2(new_n414), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(new_n408), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n416), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(new_n434), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G902), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n424), .A2(new_n415), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n452), .B2(new_n406), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n416), .A2(new_n419), .A3(new_n406), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(KEYINPUT72), .A3(new_n434), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n453), .A2(new_n447), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n443), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n441), .A2(new_n442), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(G234), .B2(new_n280), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT23), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n216), .B2(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n216), .A2(G128), .ZN(new_n463));
  INV_X1    g277(.A(new_n260), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G119), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n462), .B(new_n463), .C1(new_n465), .C2(new_n461), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G110), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT74), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT75), .B(G125), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G140), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(G125), .B2(G140), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT16), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n257), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(G146), .A3(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT24), .B(G110), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n465), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n468), .B(new_n478), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n479), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(G110), .B2(new_n466), .ZN(new_n485));
  XNOR2_X1  g299(.A(G125), .B(G140), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n257), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n477), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n402), .A2(G221), .A3(G234), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT22), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(G137), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(new_n488), .A3(new_n492), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n280), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT25), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n496), .A2(new_n498), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n460), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n495), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n492), .B1(new_n483), .B2(new_n488), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n280), .B1(new_n459), .B2(G234), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n458), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n401), .A2(new_n402), .A3(G214), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n262), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT91), .B1(new_n511), .B2(G131), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n510), .B(G143), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n412), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(G131), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n512), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(KEYINPUT17), .A3(G131), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n476), .A2(new_n477), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n521), .A2(new_n412), .A3(KEYINPUT90), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n513), .B(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n487), .B1(new_n471), .B2(new_n257), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(G113), .B(G122), .Z(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(G104), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n527), .B(KEYINPUT92), .Z(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n512), .A2(new_n517), .A3(new_n515), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT19), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n486), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n471), .B2(new_n531), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n530), .B(new_n477), .C1(G146), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n527), .B1(new_n534), .B2(new_n525), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT20), .B1(new_n538), .B2(KEYINPUT93), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n529), .B2(new_n535), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT20), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n539), .B(new_n540), .C1(new_n529), .C2(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n527), .B1(new_n520), .B2(new_n525), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n280), .B1(new_n529), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT95), .B(G475), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(G234), .A2(G237), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(G952), .A3(new_n402), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT21), .B(G898), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(G902), .A3(G953), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n262), .A2(G128), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n260), .B2(new_n262), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n321), .B1(new_n563), .B2(KEYINPUT13), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(KEYINPUT13), .B2(new_n561), .ZN(new_n565));
  INV_X1    g379(.A(G122), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G116), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(G116), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n194), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n565), .B(new_n571), .C1(G134), .C2(new_n562), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT14), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n569), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT96), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n568), .A2(KEYINPUT14), .ZN(new_n576));
  OAI21_X1  g390(.A(G107), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n194), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n562), .B(G134), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n392), .A2(new_n459), .A3(G953), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n280), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n581), .A2(new_n583), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n582), .B1(new_n572), .B2(new_n580), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n280), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n586), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n551), .A2(new_n560), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n398), .A2(new_n509), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n301), .A2(new_n599), .A3(new_n297), .A4(new_n295), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(new_n306), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n299), .A2(KEYINPUT98), .A3(new_n302), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT99), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT99), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n606), .ZN(new_n607));
  OR3_X1    g421(.A1(new_n589), .A2(new_n606), .A3(new_n590), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(new_n608), .A3(G478), .A4(new_n280), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n591), .A2(new_n585), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n551), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n605), .A2(new_n560), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n395), .A2(new_n397), .ZN(new_n615));
  INV_X1    g429(.A(new_n508), .ZN(new_n616));
  INV_X1    g430(.A(new_n440), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n443), .B1(new_n438), .B2(new_n280), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n615), .A2(KEYINPUT97), .A3(new_n616), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n601), .A2(new_n602), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT99), .ZN(new_n631));
  INV_X1    g445(.A(new_n543), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n542), .A2(KEYINPUT20), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n593), .B(new_n550), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n630), .A2(new_n560), .A3(new_n631), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n624), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT35), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n483), .A2(new_n640), .A3(new_n488), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n483), .B2(new_n488), .ZN(new_n643));
  OAI22_X1  g457(.A1(new_n642), .A2(new_n643), .B1(KEYINPUT36), .B2(new_n493), .ZN(new_n644));
  INV_X1    g458(.A(new_n643), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n641), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n506), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n496), .B(new_n498), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n460), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n398), .A2(new_n596), .A3(new_n619), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT37), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G110), .ZN(G12));
  AOI21_X1  g468(.A(new_n458), .B1(new_n395), .B2(new_n397), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n553), .B1(new_n557), .B2(G900), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n550), .B(new_n656), .C1(new_n632), .C2(new_n633), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n594), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n605), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n605), .A2(new_n655), .A3(KEYINPUT101), .A4(new_n660), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(new_n656), .B(KEYINPUT39), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n615), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n441), .A2(new_n442), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n445), .A2(new_n415), .A3(new_n434), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n280), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n452), .A2(new_n434), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n305), .B(KEYINPUT38), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n551), .A2(new_n594), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n670), .A2(new_n677), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n651), .A2(new_n307), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n681), .B(new_n682), .C1(KEYINPUT40), .C2(new_n669), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND2_X1  g498(.A1(new_n546), .A2(new_n550), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n611), .A3(new_n656), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n605), .A2(new_n655), .A3(new_n651), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(new_n375), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n374), .B1(new_n373), .B2(new_n319), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n356), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n362), .B1(new_n692), .B2(new_n345), .ZN(new_n693));
  INV_X1    g507(.A(new_n387), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n280), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n382), .A2(new_n387), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n389), .A3(new_n280), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n393), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n458), .A2(new_n699), .A3(new_n508), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n605), .A3(new_n560), .A4(new_n613), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n605), .A3(new_n560), .A4(new_n635), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  INV_X1    g519(.A(new_n699), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n458), .A2(new_n595), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n605), .A2(new_n651), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT102), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NOR2_X1   g524(.A1(new_n699), .A2(new_n680), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n427), .A2(new_n428), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n446), .A2(new_n434), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n431), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n618), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n508), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n605), .A2(new_n560), .A3(new_n711), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NOR2_X1   g532(.A1(new_n650), .A2(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n686), .A2(KEYINPUT103), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n685), .A2(new_n611), .A3(new_n721), .A4(new_n656), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n605), .A2(new_n706), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT104), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  AOI21_X1  g540(.A(new_n307), .B1(new_n303), .B2(new_n304), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n390), .A2(new_n394), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n723), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT42), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n432), .A2(new_n439), .ZN(new_n732));
  INV_X1    g546(.A(new_n457), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n508), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n728), .A3(new_n723), .A4(new_n727), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n731), .A2(new_n509), .B1(new_n735), .B2(KEYINPUT42), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n458), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n616), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n739), .A2(new_n729), .A3(new_n659), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n321), .ZN(G36));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n551), .A2(new_n611), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT43), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n650), .A2(new_n619), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT105), .Z(new_n747));
  INV_X1    g561(.A(new_n727), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n744), .A2(new_n745), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n362), .B1(new_n386), .B2(new_n345), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n692), .B2(new_n383), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n379), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n396), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n379), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n393), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n667), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n747), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  NAND2_X1  g578(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n738), .A2(new_n616), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n760), .A2(new_n767), .A3(new_n393), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n748), .A2(new_n686), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NOR2_X1   g585(.A1(new_n744), .A2(new_n553), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n716), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n765), .A2(new_n768), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n696), .A2(new_n698), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n394), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n727), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n678), .A2(new_n307), .A3(new_n706), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n773), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n748), .A2(new_n699), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n772), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT112), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n616), .A3(new_n554), .A4(new_n677), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n611), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n787), .A2(new_n719), .B1(new_n551), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n779), .B(KEYINPUT111), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT50), .B1(new_n791), .B2(new_n773), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n784), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n790), .A2(new_n792), .ZN(new_n795));
  NAND2_X1  g609(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g610(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n797));
  INV_X1    g611(.A(new_n773), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n748), .B1(new_n774), .B2(new_n776), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n605), .A3(new_n706), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n787), .A2(new_n734), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT48), .Z(new_n806));
  INV_X1    g620(.A(new_n613), .ZN(new_n807));
  OAI211_X1 g621(.A(G952), .B(new_n402), .C1(new_n788), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n593), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n588), .A2(new_n592), .A3(KEYINPUT108), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n551), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n559), .B1(new_n308), .B2(new_n310), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n622), .A2(new_n623), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n723), .A2(new_n719), .A3(new_n727), .A4(new_n728), .ZN(new_n820));
  INV_X1    g634(.A(new_n380), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n698), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT83), .B1(new_n822), .B2(new_n393), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n311), .B(new_n394), .C1(new_n698), .C2(new_n821), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n738), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n815), .A2(new_n657), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(KEYINPUT109), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n815), .A2(new_n828), .A3(new_n657), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n727), .B(new_n651), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n820), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n740), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n819), .A2(new_n832), .A3(new_n597), .A4(new_n652), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n701), .A2(new_n708), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n509), .A2(new_n706), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n636), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n630), .A2(new_n716), .A3(new_n560), .A4(new_n631), .ZN(new_n837));
  INV_X1    g651(.A(new_n711), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n840), .A3(new_n736), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n688), .A2(new_n724), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n663), .B2(new_n664), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n603), .A2(new_n604), .A3(new_n680), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n650), .A2(new_n656), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n728), .A3(new_n676), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n688), .A2(new_n724), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n665), .A2(new_n849), .A3(new_n847), .A4(KEYINPUT52), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n842), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n665), .A2(new_n849), .A3(new_n847), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n860), .B2(new_n850), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n701), .A2(new_n704), .A3(new_n708), .A4(new_n717), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n731), .A2(new_n509), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT110), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT110), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n834), .A2(new_n840), .A3(new_n867), .A4(new_n736), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n833), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n856), .A2(new_n857), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n803), .A2(new_n872), .A3(new_n804), .A4(new_n809), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n811), .A2(new_n855), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(G952), .A2(G953), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n743), .B1(new_n775), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n678), .B(new_n878), .C1(new_n877), .C2(new_n775), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n616), .A2(new_n306), .A3(new_n393), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT106), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n881), .A3(new_n676), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT107), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n280), .B1(new_n856), .B2(new_n870), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n248), .A2(new_n274), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT115), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(new_n272), .Z(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(new_n887), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n888), .A2(new_n894), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n402), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n379), .B(KEYINPUT57), .Z(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n860), .A2(new_n850), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n901), .A2(new_n869), .A3(KEYINPUT53), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n901), .B2(new_n842), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT54), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n871), .ZN(new_n905));
  INV_X1    g719(.A(new_n697), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT117), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n857), .B1(new_n856), .B2(new_n870), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n697), .ZN(new_n912));
  INV_X1    g726(.A(new_n755), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT118), .B1(new_n885), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n852), .A2(new_n853), .B1(new_n861), .B2(new_n869), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n280), .A4(new_n755), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n907), .A2(new_n912), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n897), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n536), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n897), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n855), .B2(new_n871), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n607), .A2(new_n608), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n920), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n904), .B2(new_n871), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n915), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n644), .A2(new_n647), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n897), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n504), .B(KEYINPUT119), .Z(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n915), .B2(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n939), .A2(new_n944), .A3(new_n945), .A4(new_n941), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n556), .B2(new_n270), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n819), .A2(new_n597), .A3(new_n652), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n840), .A3(new_n834), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n950), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n890), .B1(G898), .B2(new_n402), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n421), .A2(new_n423), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT121), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n533), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n402), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n817), .B(KEYINPUT123), .Z(new_n962));
  NOR4_X1   g776(.A1(new_n962), .A2(new_n739), .A3(new_n669), .A4(new_n748), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n844), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n683), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(KEYINPUT62), .A3(new_n683), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n763), .A2(new_n770), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n961), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  INV_X1    g788(.A(G900), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n360), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n740), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n845), .A2(new_n734), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n865), .B1(new_n762), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n965), .A2(new_n971), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n960), .B1(new_n980), .B2(new_n402), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n975), .A2(G953), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n973), .A2(new_n974), .A3(new_n976), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n976), .A2(new_n974), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n976), .A2(new_n974), .ZN(new_n986));
  INV_X1    g800(.A(new_n983), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n985), .B(new_n986), .C1(new_n972), .C2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n984), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(new_n968), .A2(new_n969), .ZN(new_n990));
  INV_X1    g804(.A(new_n963), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n953), .A3(new_n971), .A4(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n443), .A2(new_n280), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n674), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n451), .A2(new_n434), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n453), .A2(new_n455), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n854), .B(new_n995), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n996), .B1(new_n980), .B2(new_n952), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n434), .A3(new_n452), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1001), .A2(new_n920), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n998), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n674), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n992), .B2(new_n996), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1001), .A2(new_n920), .A3(new_n1003), .ZN(new_n1009));
  OAI21_X1  g823(.A(KEYINPUT127), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1006), .A2(new_n1010), .ZN(G57));
endmodule


