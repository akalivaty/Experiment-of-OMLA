//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT100), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n207), .B1(KEYINPUT94), .B2(new_n208), .C1(G1gat), .C2(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT94), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213));
  INV_X1    g012(.A(G64gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT99), .ZN(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G57gat), .A2(G64gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(KEYINPUT9), .ZN(new_n220));
  NAND2_X1  g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  OAI221_X1 g021(.A(new_n217), .B1(new_n215), .B2(new_n218), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n214), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n218), .C1(new_n222), .C2(KEYINPUT9), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT98), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n219), .B1(new_n226), .B2(new_n221), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n225), .B(new_n227), .C1(new_n226), .C2(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G231gat), .ZN(new_n232));
  INV_X1    g031(.A(G233gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(G231gat), .A3(G233gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n204), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(new_n213), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n241));
  INV_X1    g040(.A(G211gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n240), .B(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n237), .A3(new_n204), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n244), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n238), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G43gat), .B(G50gat), .Z(new_n251));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G29gat), .ZN(new_n254));
  INV_X1    g053(.A(G36gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT92), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT14), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(new_n254), .A3(new_n255), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n261), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT93), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(KEYINPUT15), .B2(new_n262), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n253), .A2(new_n260), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n263), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n261), .A2(KEYINPUT15), .A3(new_n262), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT17), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  INV_X1    g079(.A(G92gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(KEYINPUT8), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n280), .A2(new_n281), .B1(new_n283), .B2(KEYINPUT101), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT101), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G99gat), .B(G106gat), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n278), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G134gat), .B(G162gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n289), .ZN(new_n293));
  AND2_X1   g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n271), .A2(new_n293), .B1(KEYINPUT41), .B2(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n290), .B2(new_n295), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(KEYINPUT41), .ZN(new_n299));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n298), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n303), .B(G22gat), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(G197gat), .ZN(new_n307));
  INV_X1    g106(.A(G204gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n242), .A2(KEYINPUT77), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G211gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n313), .A3(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT22), .ZN(new_n315));
  AOI221_X4 g114(.A(G211gat), .B1(new_n309), .B2(new_n310), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n310), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n242), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n306), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT77), .B(G211gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT22), .B1(new_n321), .B2(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n318), .ZN(new_n323));
  OAI21_X1  g122(.A(G211gat), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n242), .A3(new_n318), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(G218gat), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G141gat), .B(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(G155gat), .B2(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n337));
  INV_X1    g136(.A(G141gat), .ZN(new_n338));
  INV_X1    g137(.A(G148gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n333), .A3(new_n328), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT86), .B1(new_n327), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n326), .A4(new_n320), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n344), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n320), .B2(new_n326), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT85), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n353), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  INV_X1    g162(.A(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n359), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n342), .A2(new_n333), .A3(new_n328), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n333), .B1(new_n342), .B2(new_n328), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n335), .A2(KEYINPUT80), .A3(new_n343), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n327), .A2(new_n346), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n367), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n362), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n366), .B1(new_n362), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n305), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n365), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n377), .A3(new_n366), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n304), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT3), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  INV_X1    g189(.A(G113gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT73), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G113gat), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n391), .A2(G120gat), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n388), .B(new_n389), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n389), .ZN(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(KEYINPUT1), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n387), .A2(new_n401), .A3(new_n348), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n397), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n397), .B2(new_n400), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT4), .B(new_n344), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n344), .A2(new_n400), .A3(new_n397), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n372), .A2(new_n373), .A3(new_n401), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n410), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(KEYINPUT5), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n404), .A2(new_n405), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n408), .B1(new_n417), .B2(new_n354), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n407), .A2(new_n408), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n418), .A2(new_n402), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G57gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AND4_X1   g226(.A1(KEYINPUT83), .A2(new_n422), .A3(KEYINPUT6), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n416), .B2(new_n421), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n429), .B2(KEYINPUT6), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n426), .A3(new_n421), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT82), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n416), .A2(new_n434), .A3(new_n426), .A4(new_n421), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n327), .ZN(new_n439));
  NAND2_X1  g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT24), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(G183gat), .A2(G190gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT70), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n440), .B(new_n441), .C1(KEYINPUT70), .C2(new_n443), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT25), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT23), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G169gat), .A2(G176gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n462), .A3(new_n459), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(G169gat), .B2(G176gat), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n452), .A2(new_n461), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G169gat), .ZN(new_n467));
  INV_X1    g266(.A(G176gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT23), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n465), .A3(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n469), .A2(new_n465), .A3(KEYINPUT64), .A4(new_n457), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n440), .A2(new_n443), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n446), .C1(G183gat), .C2(G190gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT25), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(KEYINPUT65), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT65), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n455), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT26), .B1(new_n481), .B2(new_n453), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n457), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n440), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G190gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT71), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT27), .B1(new_n489), .B2(new_n235), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n488), .B(new_n490), .C1(new_n491), .C2(new_n489), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G183gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT28), .A3(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT72), .B(new_n440), .C1(new_n482), .C2(new_n484), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G226gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(new_n233), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n480), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(KEYINPUT29), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n480), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n439), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n504), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n476), .A2(new_n477), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n476), .A2(KEYINPUT65), .A3(new_n477), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n462), .B1(new_n456), .B2(new_n459), .ZN(new_n512));
  INV_X1    g311(.A(new_n465), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n512), .A2(new_n451), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n510), .A2(new_n511), .B1(new_n514), .B2(new_n463), .ZN(new_n515));
  INV_X1    g314(.A(new_n499), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n507), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n480), .A2(new_n499), .A3(new_n502), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n327), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G64gat), .B(G92gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT78), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G8gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(new_n255), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n519), .A3(KEYINPUT30), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n503), .A2(new_n505), .A3(new_n439), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n327), .B1(new_n517), .B2(new_n518), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n523), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n519), .A3(KEYINPUT30), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n431), .A2(new_n438), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n386), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n418), .A2(new_n402), .A3(new_n419), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n410), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT39), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(KEYINPUT39), .C1(new_n410), .C2(new_n414), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT40), .A4(new_n426), .ZN(new_n538));
  INV_X1    g337(.A(new_n429), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n531), .A2(new_n538), .A3(new_n539), .A4(new_n524), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT40), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n537), .A3(new_n426), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n506), .A2(new_n519), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n529), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n547));
  NAND3_X1  g346(.A1(new_n506), .A2(new_n519), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT89), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n506), .A2(new_n519), .A3(new_n550), .A4(new_n547), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n549), .A2(new_n551), .B1(KEYINPUT37), .B2(new_n544), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n523), .B1(new_n552), .B2(new_n545), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n551), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n506), .A2(new_n519), .A3(KEYINPUT87), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(KEYINPUT37), .C1(KEYINPUT87), .C2(new_n519), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n546), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT6), .B(new_n429), .C1(new_n433), .C2(new_n435), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n422), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT83), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n429), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n543), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n533), .B1(new_n567), .B2(new_n386), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n570));
  INV_X1    g369(.A(new_n417), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n515), .B2(new_n516), .ZN(new_n572));
  NAND2_X1  g371(.A1(G227gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n480), .A2(new_n417), .A3(new_n499), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n572), .A2(new_n578), .A3(new_n574), .A4(new_n575), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n570), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n575), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n417), .B1(new_n480), .B2(new_n499), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n573), .B2(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI221_X1 g385(.A(new_n573), .B1(KEYINPUT76), .B2(new_n584), .C1(new_n581), .C2(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n577), .A2(new_n579), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G15gat), .B(G43gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G71gat), .B(G99gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n588), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n590), .B2(new_n591), .ZN(new_n600));
  INV_X1    g399(.A(new_n580), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n586), .A2(new_n587), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n580), .A2(new_n588), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n569), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n596), .B1(new_n589), .B2(new_n597), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n600), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT36), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n568), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n531), .A2(new_n524), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n560), .C2(new_n565), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n614), .A2(new_n385), .A3(new_n608), .A4(new_n607), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n532), .A2(new_n613), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n615), .A2(KEYINPUT35), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n385), .A2(new_n532), .A3(new_n607), .A4(new_n608), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT91), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT35), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n618), .B2(KEYINPUT35), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n250), .B(new_n302), .C1(new_n611), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n273), .A2(new_n278), .A3(new_n212), .ZN(new_n625));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  INV_X1    g426(.A(new_n212), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n271), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n271), .A2(new_n627), .A3(new_n628), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n625), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n271), .A2(new_n627), .A3(new_n628), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n633), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n637), .A2(new_n626), .A3(new_n625), .A4(new_n638), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n630), .A2(new_n629), .B1(new_n271), .B2(new_n628), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n626), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT11), .B(G169gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G197gat), .ZN(new_n646));
  XOR2_X1   g445(.A(G113gat), .B(G141gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n639), .A3(new_n649), .A4(new_n643), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n289), .A2(new_n229), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n289), .A2(new_n229), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n289), .A2(new_n229), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT10), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G230gat), .ZN(new_n662));
  OAI22_X1  g461(.A1(new_n659), .A2(new_n661), .B1(new_n662), .B2(new_n233), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n233), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n656), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT103), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G120gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n339), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n671), .A2(KEYINPUT104), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT104), .B1(new_n671), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n653), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n624), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n566), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n679), .A2(new_n612), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n612), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n208), .B1(new_n680), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n685), .A2(KEYINPUT105), .A3(KEYINPUT42), .A4(new_n686), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(G1325gat));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT36), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT36), .B1(new_n607), .B2(new_n608), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n606), .A2(KEYINPUT106), .A3(new_n609), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n680), .A2(G15gat), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n598), .A2(new_n605), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n680), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n679), .A2(new_n385), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n568), .A2(new_n700), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n623), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n302), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n302), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n611), .B2(new_n623), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n250), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(new_n653), .A3(new_n677), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n566), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n717), .A2(new_n722), .A3(new_n566), .A4(new_n719), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(G29gat), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n715), .A2(new_n719), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n254), .A3(new_n566), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n255), .A3(new_n690), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n717), .A2(new_n690), .A3(new_n719), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n255), .ZN(G1329gat));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n716), .A3(G43gat), .A4(new_n719), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(new_n700), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n703), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n725), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n736), .A2(new_n737), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n735), .B2(new_n700), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n740), .B(new_n741), .C1(new_n735), .C2(new_n700), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n744), .A3(new_n746), .ZN(G1330gat));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n716), .A3(new_n386), .A4(new_n719), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G50gat), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT48), .B1(new_n749), .B2(KEYINPUT111), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n386), .A2(new_n364), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT110), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n751), .A2(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n749), .B(new_n754), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1331gat));
  INV_X1    g557(.A(new_n653), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n709), .B2(new_n623), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n250), .A2(new_n676), .A3(new_n302), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n566), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n216), .ZN(G1332gat));
  NAND2_X1  g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n760), .A2(new_n690), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n768), .B(new_n769), .Z(G1333gat));
  NAND4_X1  g569(.A1(new_n760), .A2(G71gat), .A3(new_n701), .A4(new_n761), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n762), .A2(new_n739), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G71gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g573(.A1(new_n762), .A2(new_n385), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g575(.A1(new_n250), .A2(new_n653), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT113), .Z(new_n778));
  NAND4_X1  g577(.A1(new_n713), .A2(new_n716), .A3(new_n677), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n763), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n557), .B(new_n523), .C1(new_n545), .C2(new_n552), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n763), .B1(new_n781), .B2(new_n546), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n385), .B1(new_n782), .B2(new_n543), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n783), .A2(new_n533), .B1(new_n698), .B2(new_n699), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n615), .A2(KEYINPUT35), .A3(new_n616), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT91), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n620), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n302), .B(new_n778), .C1(new_n784), .C2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n302), .A4(new_n778), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n280), .B(new_n677), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n780), .B1(new_n796), .B2(new_n763), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n779), .B2(new_n612), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n791), .A2(new_n793), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n281), .A3(new_n677), .A4(new_n690), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n739), .A2(G99gat), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n677), .B(new_n806), .C1(new_n794), .C2(new_n795), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n779), .B2(new_n700), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  OAI21_X1  g612(.A(G106gat), .B1(new_n779), .B2(new_n385), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n385), .A2(new_n676), .A3(G106gat), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n763), .A2(new_n690), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n626), .B1(new_n637), .B2(new_n625), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n640), .A2(new_n642), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n648), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n652), .B(new_n826), .C1(new_n674), .C2(new_n675), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n659), .A2(new_n661), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n664), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(KEYINPUT54), .A3(new_n663), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n663), .A2(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n670), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT55), .A4(new_n670), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n673), .A3(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n714), .B(new_n827), .C1(new_n653), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n652), .A2(new_n826), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n302), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n250), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n718), .A2(new_n653), .A3(new_n676), .A4(new_n714), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n386), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  AOI211_X1 g643(.A(new_n844), .B(new_n386), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n703), .B(new_n823), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n653), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n842), .A2(new_n566), .A3(new_n703), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n690), .B1(new_n848), .B2(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n392), .A2(new_n394), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n847), .B1(new_n855), .B2(new_n653), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n846), .B2(new_n676), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n677), .A2(new_n390), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n861), .A3(new_n250), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n849), .A2(new_n718), .A3(new_n850), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(G1342gat));
  NOR3_X1   g663(.A1(new_n851), .A2(G134gat), .A3(new_n714), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n846), .B2(new_n714), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n385), .B1(new_n840), .B2(new_n841), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT57), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n700), .A3(new_n823), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n653), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n840), .A2(new_n841), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n386), .A2(new_n875), .A3(new_n700), .A4(new_n823), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n338), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n653), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n339), .A3(new_n677), .ZN(new_n880));
  INV_X1    g679(.A(new_n873), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n677), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(G148gat), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n882), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(G155gat), .B1(new_n876), .B2(new_n718), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n718), .A2(G155gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT120), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n881), .B2(new_n890), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n892), .A3(new_n302), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT121), .ZN(new_n894));
  OAI21_X1  g693(.A(G162gat), .B1(new_n873), .B2(new_n714), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n875), .A2(new_n763), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT122), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n899), .A3(new_n763), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n739), .A2(new_n386), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(new_n690), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n467), .A3(new_n759), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n566), .A2(new_n612), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n703), .B(new_n905), .C1(new_n843), .C2(new_n845), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n653), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(G1348gat));
  NOR3_X1   g707(.A1(new_n906), .A2(new_n468), .A3(new_n676), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n903), .A2(new_n677), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n468), .ZN(G1349gat));
  OAI21_X1  g710(.A(G183gat), .B1(new_n906), .B2(new_n250), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n718), .A2(new_n495), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n901), .A2(new_n690), .A3(new_n902), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(KEYINPUT123), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(KEYINPUT123), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n912), .A2(new_n915), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n919), .B2(new_n922), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n903), .A2(new_n488), .A3(new_n302), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n906), .A2(new_n714), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(G190gat), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n925), .B2(G190gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n872), .A2(new_n700), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n931), .A2(KEYINPUT126), .A3(new_n759), .A4(new_n905), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n872), .A2(new_n700), .A3(new_n905), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n653), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(G197gat), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n701), .A2(new_n385), .A3(new_n612), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n901), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n307), .A3(new_n759), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n941), .ZN(G1352gat));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n308), .A3(new_n677), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n934), .A2(KEYINPUT127), .A3(new_n676), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(new_n934), .B2(new_n676), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(G204gat), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(G1353gat));
  INV_X1    g748(.A(new_n321), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n940), .A2(new_n950), .A3(new_n718), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n718), .A3(new_n905), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n306), .A3(new_n302), .ZN(new_n957));
  OAI21_X1  g756(.A(G218gat), .B1(new_n934), .B2(new_n714), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


