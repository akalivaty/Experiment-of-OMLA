//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT81), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G106gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT71), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT74), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G141gat), .B(G148gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n224), .B2(new_n225), .ZN(new_n228));
  OAI221_X1 g027(.A(new_n217), .B1(new_n220), .B2(new_n223), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT76), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n217), .B1(new_n221), .B2(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT77), .B(G141gat), .ZN(new_n232));
  INV_X1    g031(.A(G148gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G141gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(G148gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n231), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n216), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n212), .A2(new_n240), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n230), .A2(new_n237), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(KEYINPUT80), .B(new_n245), .C1(new_n241), .C2(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT3), .B1(new_n216), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n237), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n256), .A2(new_n245), .A3(new_n241), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n251), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G78gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT80), .B1(new_n244), .B2(new_n245), .ZN(new_n260));
  INV_X1    g059(.A(new_n249), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G22gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n259), .B1(new_n258), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n205), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n251), .B1(new_n250), .B2(new_n257), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n262), .A2(G22gat), .ZN(new_n269));
  OAI21_X1  g068(.A(G78gat), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n264), .A3(new_n204), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT26), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n276), .B(KEYINPUT66), .Z(new_n280));
  OAI211_X1 g079(.A(new_n278), .B(new_n279), .C1(KEYINPUT26), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n283), .B2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n284), .A2(new_n285), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n281), .B(new_n286), .C1(new_n285), .C2(new_n284), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(new_n274), .C1(KEYINPUT23), .C2(new_n276), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT64), .Z(new_n293));
  NOR2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT25), .B1(new_n280), .B2(new_n295), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n294), .A2(KEYINPUT25), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT1), .ZN(new_n300));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n300), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G227gat), .A2(G233gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n304), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT34), .B1(new_n309), .B2(KEYINPUT70), .ZN(new_n310));
  XOR2_X1   g109(.A(G15gat), .B(G43gat), .Z(new_n311));
  XNOR2_X1  g110(.A(G71gat), .B(G99gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(KEYINPUT33), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n315), .A2(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(new_n310), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n298), .B2(new_n252), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n298), .A2(new_n336), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n215), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n298), .ZN(new_n344));
  INV_X1    g143(.A(new_n240), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n216), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n334), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n339), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n342), .B1(new_n337), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n216), .ZN(new_n351));
  INV_X1    g150(.A(new_n347), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n333), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(KEYINPUT30), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n343), .A2(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n333), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n267), .A2(new_n271), .A3(new_n330), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n255), .A2(new_n304), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n254), .A2(new_n305), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n305), .A3(new_n239), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n371), .A2(new_n373), .A3(new_n374), .A4(new_n365), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT79), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n370), .B1(new_n375), .B2(KEYINPUT79), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n364), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(KEYINPUT79), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT5), .A3(new_n369), .ZN(new_n381));
  INV_X1    g180(.A(new_n364), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n376), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT82), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT35), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n360), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n387), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT35), .B1(new_n359), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT36), .ZN(new_n395));
  INV_X1    g194(.A(new_n329), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n326), .B1(new_n321), .B2(new_n324), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n328), .A2(KEYINPUT36), .A3(new_n329), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n267), .A2(new_n271), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n387), .A2(new_n358), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n265), .A2(new_n266), .A3(new_n205), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n204), .B1(new_n270), .B2(new_n264), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT38), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n333), .B1(new_n355), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n351), .A2(new_n352), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT37), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n350), .A2(new_n215), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n346), .A2(new_n340), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n414), .B2(new_n216), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT38), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(new_n334), .C1(KEYINPUT37), .C2(new_n410), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n353), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n388), .A2(new_n419), .A3(new_n390), .ZN(new_n420));
  INV_X1    g219(.A(new_n358), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n366), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT39), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n367), .A2(new_n368), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n423), .B(KEYINPUT39), .C1(new_n366), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n426), .A3(new_n364), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT40), .A4(new_n364), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n421), .A2(new_n383), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n420), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n392), .A2(new_n394), .B1(new_n403), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n436));
  INV_X1    g235(.A(G29gat), .ZN(new_n437));
  INV_X1    g236(.A(G36gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G29gat), .A2(G36gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n435), .A2(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(G43gat), .A2(G50gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(G43gat), .A2(G50gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT15), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n451), .B(KEYINPUT85), .C1(new_n448), .C2(new_n444), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459));
  INV_X1    g258(.A(G1gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT16), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n459), .A2(G1gat), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(G8gat), .ZN(new_n464));
  INV_X1    g263(.A(G8gat), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n459), .A2(G1gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n461), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(G8gat), .B1(new_n462), .B2(new_n463), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n465), .A3(new_n467), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT86), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT86), .B1(new_n470), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT87), .B1(new_n474), .B2(new_n454), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n464), .B2(new_n468), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT86), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n452), .A2(new_n453), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n458), .A2(new_n469), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT18), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n455), .A2(new_n469), .A3(new_n457), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n454), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n479), .B2(new_n480), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT18), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT88), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n475), .A2(new_n482), .B1(new_n454), .B2(new_n474), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n485), .B(KEYINPUT13), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n474), .A2(new_n454), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n488), .B2(new_n489), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n494), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n434), .B1(new_n493), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G197gat), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT11), .B(G169gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n508), .B(KEYINPUT12), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n434), .B(new_n511), .C1(new_n493), .C2(new_n503), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n433), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G99gat), .B(G106gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g316(.A(G92gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G92gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G99gat), .ZN(new_n524));
  INV_X1    g323(.A(G106gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT8), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT92), .B1(new_n523), .B2(new_n526), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n515), .B(new_n517), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n515), .B1(new_n535), .B2(new_n517), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n458), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n480), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G190gat), .B(G218gat), .Z(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  XOR2_X1   g342(.A(G134gat), .B(G162gat), .Z(new_n544));
  AOI21_X1  g343(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n546), .B(KEYINPUT93), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G71gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n259), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n555), .A2(KEYINPUT90), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G127gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n479), .B1(KEYINPUT21), .B2(new_n559), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G155gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n566), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT94), .ZN(new_n573));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n556), .B(new_n558), .Z(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n536), .B2(new_n530), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n517), .B1(new_n527), .B2(new_n528), .ZN(new_n578));
  INV_X1    g377(.A(new_n515), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n559), .A3(new_n529), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n538), .A2(KEYINPUT95), .A3(new_n559), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT10), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n580), .A2(new_n559), .A3(KEYINPUT10), .A4(new_n529), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n574), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(KEYINPUT97), .B(new_n574), .C1(new_n584), .C2(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(new_n574), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n592), .A3(new_n583), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  AND2_X1   g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT98), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n590), .A2(new_n600), .A3(new_n591), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n588), .A2(new_n593), .ZN(new_n603));
  INV_X1    g402(.A(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n573), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n514), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n387), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n460), .ZN(G1324gat));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n358), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(KEYINPUT100), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(KEYINPUT100), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(G8gat), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(KEYINPUT42), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(KEYINPUT101), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n620));
  OAI211_X1 g419(.A(new_n615), .B(new_n617), .C1(new_n619), .C2(new_n620), .ZN(G1325gat));
  AND2_X1   g420(.A1(new_n398), .A2(new_n399), .ZN(new_n622));
  OAI21_X1  g421(.A(G15gat), .B1(new_n609), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n330), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n624), .A2(G15gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n609), .B2(new_n625), .ZN(G1326gat));
  NOR3_X1   g425(.A1(new_n433), .A2(new_n406), .A3(new_n513), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n608), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  NOR3_X1   g429(.A1(new_n551), .A2(new_n571), .A3(new_n606), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n514), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n632), .A2(G29gat), .A3(new_n387), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT45), .Z(new_n634));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n433), .B2(new_n551), .ZN(new_n636));
  INV_X1    g435(.A(new_n551), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n406), .A2(new_n387), .A3(new_n358), .A4(new_n330), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n638), .A2(KEYINPUT35), .B1(new_n360), .B2(new_n391), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n640));
  INV_X1    g439(.A(new_n390), .ZN(new_n641));
  NOR4_X1   g440(.A1(new_n640), .A2(new_n641), .A3(new_n412), .A4(new_n418), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n431), .A2(new_n267), .A3(new_n271), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT44), .B(new_n637), .C1(new_n639), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n636), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n513), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n571), .B(KEYINPUT103), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n649), .A2(new_n607), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n387), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n634), .A2(new_n654), .ZN(G1328gat));
  NOR3_X1   g454(.A1(new_n632), .A2(G36gat), .A3(new_n358), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT46), .ZN(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n653), .B2(new_n358), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1329gat));
  OAI21_X1  g458(.A(G43gat), .B1(new_n653), .B2(new_n622), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n632), .A2(G43gat), .A3(new_n624), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n660), .B2(new_n662), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(G1330gat));
  OAI21_X1  g464(.A(G50gat), .B1(new_n653), .B2(new_n406), .ZN(new_n666));
  INV_X1    g465(.A(G50gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n627), .A2(new_n667), .A3(new_n631), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT48), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(KEYINPUT48), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1331gat));
  NAND2_X1  g472(.A1(new_n392), .A2(new_n394), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n403), .A2(new_n432), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n651), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n573), .A2(new_n677), .A3(new_n606), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n387), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT104), .B(G57gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1332gat));
  NOR2_X1   g481(.A1(new_n679), .A2(new_n358), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n684));
  AND2_X1   g483(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n683), .B2(new_n684), .ZN(G1333gat));
  NAND4_X1  g486(.A1(new_n676), .A2(G71gat), .A3(new_n400), .A4(new_n678), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT105), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n552), .B1(new_n679), .B2(new_n624), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1334gat));
  NOR2_X1   g492(.A1(new_n679), .A2(new_n406), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n259), .ZN(G1335gat));
  NOR3_X1   g494(.A1(new_n651), .A2(new_n571), .A3(new_n607), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n649), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G85gat), .B1(new_n698), .B2(new_n387), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n433), .A2(new_n551), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n651), .A2(new_n571), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT51), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND4_X1   g501(.A1(KEYINPUT51), .A2(new_n676), .A3(new_n637), .A4(new_n701), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n606), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n393), .A2(new_n522), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n699), .B1(new_n705), .B2(new_n706), .ZN(G1336gat));
  NOR2_X1   g506(.A1(new_n358), .A2(G92gat), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n606), .B(new_n708), .C1(new_n702), .C2(new_n703), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n636), .A2(new_n648), .A3(new_n421), .A4(new_n697), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n519), .A2(new_n521), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n709), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n712), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n709), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT52), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n718), .B2(KEYINPUT52), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n714), .B1(new_n720), .B2(new_n721), .ZN(G1337gat));
  NOR3_X1   g521(.A1(new_n698), .A2(new_n524), .A3(new_n622), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n330), .A3(new_n606), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n524), .ZN(G1338gat));
  OAI21_X1  g524(.A(G106gat), .B1(new_n698), .B2(new_n406), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n401), .A2(new_n525), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n705), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g528(.A(KEYINPUT54), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n582), .A2(new_n583), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT10), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n585), .A2(KEYINPUT96), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n585), .A2(KEYINPUT96), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n731), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n730), .B1(new_n735), .B2(new_n592), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n590), .A3(new_n591), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n738));
  OAI211_X1 g537(.A(new_n574), .B(new_n738), .C1(new_n584), .C2(new_n587), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n604), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n740), .A3(KEYINPUT55), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n602), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n602), .A2(KEYINPUT111), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n737), .A2(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n651), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n483), .A2(new_n485), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n501), .A2(new_n496), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n508), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n493), .A2(new_n503), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n511), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n606), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n637), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n753), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n551), .A2(new_n758), .ZN(new_n759));
  AND4_X1   g558(.A1(new_n745), .A2(new_n759), .A3(new_n748), .A4(new_n744), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n652), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n608), .A2(new_n677), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n387), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n360), .ZN(new_n764));
  INV_X1    g563(.A(G113gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n513), .ZN(new_n766));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n651), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n765), .B2(new_n768), .ZN(G1340gat));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n606), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G120gat), .ZN(G1341gat));
  NOR3_X1   g570(.A1(new_n764), .A2(new_n563), .A3(new_n652), .ZN(new_n772));
  INV_X1    g571(.A(new_n571), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(G127gat), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT112), .B1(new_n764), .B2(new_n773), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1342gat));
  NOR2_X1   g576(.A1(new_n421), .A2(new_n551), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n763), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n401), .A2(new_n624), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(G134gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n786), .A3(new_n782), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT114), .Z(new_n789));
  AOI21_X1  g588(.A(new_n785), .B1(new_n784), .B2(new_n787), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n780), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(G134gat), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1343gat));
  NOR3_X1   g592(.A1(new_n400), .A2(new_n387), .A3(new_n421), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n406), .B1(new_n761), .B2(new_n762), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(KEYINPUT57), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n401), .A2(KEYINPUT57), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n748), .A2(KEYINPUT115), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n746), .A2(new_n799), .A3(new_n747), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n510), .A2(new_n602), .A3(new_n512), .A4(new_n741), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n756), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT116), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n756), .B(new_n805), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n551), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n760), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n571), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n797), .B1(new_n810), .B2(new_n762), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n794), .B1(new_n796), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n232), .B1(new_n812), .B2(new_n513), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n795), .A2(new_n393), .A3(new_n622), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n358), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n510), .A2(new_n235), .A3(new_n512), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n813), .B(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n812), .A2(new_n677), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n232), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n814), .ZN(G1344gat));
  NOR2_X1   g621(.A1(new_n233), .A2(KEYINPUT59), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n812), .B2(new_n607), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n797), .B1(new_n761), .B2(new_n762), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n573), .A2(new_n513), .A3(new_n607), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT118), .B1(new_n809), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n637), .B1(new_n803), .B2(KEYINPUT116), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n760), .B1(new_n830), .B2(new_n806), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n829), .B(new_n826), .C1(new_n831), .C2(new_n571), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n401), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n825), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n794), .A2(new_n606), .ZN(new_n836));
  OAI21_X1  g635(.A(G148gat), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n824), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n606), .A2(new_n233), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n816), .B2(new_n843), .ZN(G1345gat));
  NOR3_X1   g643(.A1(new_n812), .A2(new_n218), .A3(new_n652), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n816), .A2(KEYINPUT120), .A3(new_n773), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(G155gat), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n816), .B2(new_n773), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G1346gat));
  OAI21_X1  g648(.A(G162gat), .B1(new_n812), .B2(new_n551), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n815), .A2(new_n219), .A3(new_n778), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1347gat));
  AOI21_X1  g651(.A(new_n393), .B1(new_n761), .B2(new_n762), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n781), .A2(new_n358), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(G169gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(new_n513), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n853), .B(KEYINPUT121), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n651), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n860), .B2(new_n856), .ZN(G1348gat));
  INV_X1    g660(.A(G176gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n606), .ZN(new_n863));
  OAI21_X1  g662(.A(G176gat), .B1(new_n855), .B2(new_n607), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1349gat));
  NAND3_X1  g664(.A1(new_n859), .A2(new_n282), .A3(new_n571), .ZN(new_n866));
  OAI21_X1  g665(.A(G183gat), .B1(new_n855), .B2(new_n652), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1350gat));
  INV_X1    g669(.A(G190gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n859), .A2(new_n871), .A3(new_n637), .ZN(new_n872));
  OAI21_X1  g671(.A(G190gat), .B1(new_n855), .B2(new_n551), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT61), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1351gat));
  NOR2_X1   g674(.A1(new_n400), .A2(new_n358), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n393), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n835), .B2(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n826), .B1(new_n831), .B2(new_n571), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n406), .B1(new_n882), .B2(KEYINPUT118), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n883), .B2(new_n832), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(new_n825), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(G197gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n513), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n877), .A2(new_n406), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n858), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(G197gat), .B1(new_n890), .B2(new_n651), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(G1352gat));
  XNOR2_X1  g691(.A(KEYINPUT124), .B(G204gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n607), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n858), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT62), .Z(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n886), .B2(new_n607), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n207), .A3(new_n571), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n571), .ZN(new_n900));
  OAI21_X1  g699(.A(G211gat), .B1(new_n835), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(G1354gat));
  NAND3_X1  g705(.A1(new_n858), .A2(new_n637), .A3(new_n889), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n208), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n833), .A2(new_n834), .ZN(new_n909));
  INV_X1    g708(.A(new_n825), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(KEYINPUT123), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n885), .A2(new_n911), .A3(KEYINPUT125), .A4(new_n878), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n551), .A2(new_n208), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT126), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT125), .B1(new_n880), .B2(new_n885), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT127), .B(new_n908), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1355gat));
endmodule


