

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U553 ( .A(n888), .Z(n520) );
  NOR2_X1 U554 ( .A1(G2104), .A2(n525), .ZN(n888) );
  NOR2_X2 U555 ( .A1(n526), .A2(n525), .ZN(n887) );
  OR2_X1 U556 ( .A1(n658), .A2(n652), .ZN(n657) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n675) );
  INV_X1 U558 ( .A(KEYINPUT103), .ZN(n699) );
  XNOR2_X1 U559 ( .A(n700), .B(n699), .ZN(n706) );
  XNOR2_X1 U560 ( .A(n708), .B(KEYINPUT32), .ZN(n735) );
  AND2_X1 U561 ( .A1(n735), .A2(n719), .ZN(n726) );
  INV_X1 U562 ( .A(KEYINPUT71), .ZN(n636) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n628) );
  INV_X1 U564 ( .A(KEYINPUT65), .ZN(n609) );
  XOR2_X1 U565 ( .A(KEYINPUT15), .B(n640), .Z(n865) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n797) );
  XNOR2_X1 U567 ( .A(KEYINPUT87), .B(n532), .ZN(G164) );
  INV_X1 U568 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2105), .A2(n526), .ZN(n604) );
  BUF_X1 U570 ( .A(n604), .Z(n892) );
  NAND2_X1 U571 ( .A1(n892), .A2(G102), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n521), .B(KEYINPUT86), .ZN(n531) );
  INV_X1 U573 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U574 ( .A1(G126), .A2(n520), .ZN(n524) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n522), .Z(n601) );
  NAND2_X1 U577 ( .A1(G138), .A2(n601), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G114), .A2(n887), .ZN(n527) );
  XNOR2_X1 U580 ( .A(KEYINPUT85), .B(n527), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n566) );
  NOR2_X2 U584 ( .A1(G651), .A2(n566), .ZN(n800) );
  NAND2_X1 U585 ( .A1(G52), .A2(n800), .ZN(n535) );
  INV_X1 U586 ( .A(G651), .ZN(n536) );
  NOR2_X1 U587 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n533), .Z(n801) );
  NAND2_X1 U589 ( .A1(G64), .A2(n801), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X2 U591 ( .A1(n566), .A2(n536), .ZN(n796) );
  NAND2_X1 U592 ( .A1(G77), .A2(n796), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G90), .A2(n797), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT67), .B(n542), .Z(G171) );
  INV_X1 U598 ( .A(G171), .ZN(G301) );
  XOR2_X1 U599 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n543) );
  XNOR2_X1 U600 ( .A(KEYINPUT5), .B(n543), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G89), .A2(n797), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n544), .B(KEYINPUT72), .ZN(n545) );
  XNOR2_X1 U603 ( .A(n545), .B(KEYINPUT4), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G76), .A2(n796), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n549), .B(n548), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G51), .A2(n800), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G63), .A2(n801), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G75), .A2(n796), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G88), .A2(n797), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G50), .A2(n800), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G62), .A2(n801), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(G166) );
  INV_X1 U621 ( .A(G166), .ZN(G303) );
  NAND2_X1 U622 ( .A1(G49), .A2(n800), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G74), .A2(G651), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U625 ( .A(KEYINPUT80), .B(n564), .ZN(n565) );
  NOR2_X1 U626 ( .A1(n801), .A2(n565), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n566), .A2(G87), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G288) );
  NAND2_X1 U629 ( .A1(G73), .A2(n796), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT2), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G86), .A2(n797), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G61), .A2(n801), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G48), .A2(n800), .ZN(n572) );
  XNOR2_X1 U635 ( .A(KEYINPUT81), .B(n572), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(G305) );
  NAND2_X1 U638 ( .A1(G72), .A2(n796), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G85), .A2(n797), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G60), .A2(n801), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT66), .B(n579), .Z(n580) );
  NOR2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n800), .A2(G47), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U646 ( .A1(G129), .A2(n520), .ZN(n585) );
  BUF_X1 U647 ( .A(n601), .Z(n895) );
  NAND2_X1 U648 ( .A1(G141), .A2(n895), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G105), .A2(n892), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT38), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT93), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n887), .A2(G117), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n909) );
  AND2_X1 U656 ( .A1(n909), .A2(G1996), .ZN(n934) );
  NAND2_X1 U657 ( .A1(G95), .A2(n892), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G131), .A2(n895), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n594), .B(KEYINPUT91), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G107), .A2(n887), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n520), .A2(G119), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT90), .B(n597), .Z(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT92), .B(n600), .Z(n900) );
  AND2_X1 U667 ( .A1(G1991), .A2(n900), .ZN(n946) );
  OR2_X1 U668 ( .A1(n934), .A2(n946), .ZN(n614) );
  NAND2_X1 U669 ( .A1(G113), .A2(n887), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G137), .A2(n601), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n612) );
  NAND2_X1 U672 ( .A1(n888), .A2(G125), .ZN(n608) );
  NAND2_X1 U673 ( .A1(n604), .A2(G101), .ZN(n606) );
  INV_X1 U674 ( .A(KEYINPUT23), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U679 ( .A(KEYINPUT64), .B(n613), .ZN(G160) );
  NAND2_X1 U680 ( .A1(G40), .A2(G160), .ZN(n626) );
  NOR2_X1 U681 ( .A1(n628), .A2(n626), .ZN(n765) );
  NAND2_X1 U682 ( .A1(n614), .A2(n765), .ZN(n752) );
  XNOR2_X1 U683 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G116), .A2(n887), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G128), .A2(n520), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT35), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n624) );
  NAND2_X1 U689 ( .A1(G104), .A2(n892), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G140), .A2(n895), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U692 ( .A(KEYINPUT34), .B(n622), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U694 ( .A(KEYINPUT36), .B(n625), .ZN(n904) );
  XNOR2_X1 U695 ( .A(KEYINPUT37), .B(G2067), .ZN(n763) );
  NOR2_X1 U696 ( .A1(n904), .A2(n763), .ZN(n954) );
  NAND2_X1 U697 ( .A1(n765), .A2(n954), .ZN(n760) );
  NAND2_X1 U698 ( .A1(n752), .A2(n760), .ZN(n749) );
  INV_X1 U699 ( .A(n626), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n687) );
  INV_X1 U701 ( .A(n687), .ZN(n682) );
  AND2_X1 U702 ( .A1(n682), .A2(G1996), .ZN(n629) );
  XOR2_X1 U703 ( .A(n629), .B(KEYINPUT26), .Z(n631) );
  INV_X1 U704 ( .A(n682), .ZN(n701) );
  NAND2_X1 U705 ( .A1(n701), .A2(G1341), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n658) );
  NAND2_X1 U707 ( .A1(G92), .A2(n797), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G66), .A2(n801), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n639) );
  NAND2_X1 U710 ( .A1(G79), .A2(n796), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G54), .A2(n800), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  INV_X1 U715 ( .A(n865), .ZN(n651) );
  NAND2_X1 U716 ( .A1(G56), .A2(n801), .ZN(n641) );
  XOR2_X1 U717 ( .A(KEYINPUT14), .B(n641), .Z(n648) );
  NAND2_X1 U718 ( .A1(G81), .A2(n797), .ZN(n642) );
  XOR2_X1 U719 ( .A(KEYINPUT12), .B(n642), .Z(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT69), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G68), .A2(n796), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT13), .B(n646), .Z(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n800), .A2(G43), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n986) );
  OR2_X1 U727 ( .A1(n651), .A2(n986), .ZN(n652) );
  XOR2_X1 U728 ( .A(KEYINPUT97), .B(n687), .Z(n680) );
  INV_X1 U729 ( .A(n680), .ZN(n662) );
  NAND2_X1 U730 ( .A1(G2067), .A2(n662), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G1348), .A2(n701), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U733 ( .A(KEYINPUT100), .B(n655), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n986), .A2(n658), .ZN(n659) );
  OR2_X1 U736 ( .A1(n865), .A2(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n662), .A2(G2072), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT27), .ZN(n665) );
  XNOR2_X1 U740 ( .A(G1956), .B(KEYINPUT99), .ZN(n1013) );
  NOR2_X1 U741 ( .A1(n1013), .A2(n662), .ZN(n664) );
  NOR2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n674) );
  NAND2_X1 U743 ( .A1(G53), .A2(n800), .ZN(n667) );
  NAND2_X1 U744 ( .A1(G65), .A2(n801), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G78), .A2(n796), .ZN(n669) );
  NAND2_X1 U747 ( .A1(G91), .A2(n797), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n929) );
  NAND2_X1 U750 ( .A1(n674), .A2(n929), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n678) );
  NOR2_X1 U752 ( .A1(n674), .A2(n929), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(KEYINPUT29), .ZN(n686) );
  XOR2_X1 U756 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NOR2_X1 U757 ( .A1(n961), .A2(n680), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(KEYINPUT98), .ZN(n684) );
  XNOR2_X1 U759 ( .A(G1961), .B(KEYINPUT96), .ZN(n1005) );
  NOR2_X1 U760 ( .A1(n1005), .A2(n682), .ZN(n683) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n692) );
  NOR2_X1 U762 ( .A1(G301), .A2(n692), .ZN(n685) );
  NOR2_X1 U763 ( .A1(n686), .A2(n685), .ZN(n697) );
  NAND2_X1 U764 ( .A1(G8), .A2(n701), .ZN(n743) );
  NOR2_X1 U765 ( .A1(G1966), .A2(n743), .ZN(n711) );
  NOR2_X1 U766 ( .A1(n687), .A2(G2084), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n713), .B(KEYINPUT95), .ZN(n688) );
  NAND2_X1 U768 ( .A1(G8), .A2(n688), .ZN(n689) );
  NOR2_X1 U769 ( .A1(n711), .A2(n689), .ZN(n690) );
  XOR2_X1 U770 ( .A(KEYINPUT30), .B(n690), .Z(n691) );
  NOR2_X1 U771 ( .A1(G168), .A2(n691), .ZN(n694) );
  AND2_X1 U772 ( .A1(G301), .A2(n692), .ZN(n693) );
  NOR2_X1 U773 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U774 ( .A(n695), .B(KEYINPUT31), .ZN(n696) );
  NOR2_X1 U775 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U776 ( .A(n698), .B(KEYINPUT101), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n709), .A2(G286), .ZN(n700) );
  NOR2_X1 U778 ( .A1(G1971), .A2(n743), .ZN(n703) );
  NOR2_X1 U779 ( .A1(G2090), .A2(n701), .ZN(n702) );
  NOR2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U781 ( .A1(G303), .A2(n704), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U783 ( .A1(n707), .A2(G8), .ZN(n708) );
  INV_X1 U784 ( .A(n709), .ZN(n710) );
  NOR2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U786 ( .A(KEYINPUT102), .B(n712), .ZN(n716) );
  XOR2_X1 U787 ( .A(KEYINPUT95), .B(n713), .Z(n714) );
  NAND2_X1 U788 ( .A1(G8), .A2(n714), .ZN(n715) );
  NAND2_X1 U789 ( .A1(n716), .A2(n715), .ZN(n734) );
  NAND2_X1 U790 ( .A1(G1976), .A2(G288), .ZN(n983) );
  INV_X1 U791 ( .A(n743), .ZN(n717) );
  NAND2_X1 U792 ( .A1(n983), .A2(n717), .ZN(n722) );
  INV_X1 U793 ( .A(n722), .ZN(n718) );
  AND2_X1 U794 ( .A1(n734), .A2(n718), .ZN(n719) );
  NOR2_X1 U795 ( .A1(G1976), .A2(G288), .ZN(n728) );
  NOR2_X1 U796 ( .A1(G1971), .A2(G303), .ZN(n720) );
  NOR2_X1 U797 ( .A1(n728), .A2(n720), .ZN(n992) );
  XNOR2_X1 U798 ( .A(KEYINPUT104), .B(n992), .ZN(n721) );
  OR2_X1 U799 ( .A1(n722), .A2(n721), .ZN(n724) );
  INV_X1 U800 ( .A(KEYINPUT33), .ZN(n723) );
  NAND2_X1 U801 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n733) );
  XNOR2_X1 U803 ( .A(G1981), .B(KEYINPUT105), .ZN(n727) );
  XNOR2_X1 U804 ( .A(n727), .B(G305), .ZN(n993) );
  INV_X1 U805 ( .A(n993), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n728), .A2(KEYINPUT33), .ZN(n729) );
  NOR2_X1 U807 ( .A1(n743), .A2(n729), .ZN(n730) );
  OR2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n747) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U811 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U812 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n739), .A2(n743), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1981), .A2(G305), .ZN(n740) );
  XOR2_X1 U816 ( .A(n740), .B(KEYINPUT24), .Z(n741) );
  XNOR2_X1 U817 ( .A(KEYINPUT94), .B(n741), .ZN(n742) );
  OR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U823 ( .A1(n990), .A2(n765), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n768) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n909), .ZN(n943) );
  INV_X1 U826 ( .A(n752), .ZN(n756) );
  NOR2_X1 U827 ( .A1(G1991), .A2(n900), .ZN(n933) );
  NOR2_X1 U828 ( .A1(G1986), .A2(G290), .ZN(n753) );
  XNOR2_X1 U829 ( .A(KEYINPUT106), .B(n753), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n933), .A2(n754), .ZN(n755) );
  NOR2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U832 ( .A1(n943), .A2(n757), .ZN(n759) );
  XOR2_X1 U833 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n758) );
  XNOR2_X1 U834 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n762), .B(KEYINPUT108), .ZN(n764) );
  NAND2_X1 U837 ( .A1(n904), .A2(n763), .ZN(n951) );
  NAND2_X1 U838 ( .A1(n764), .A2(n951), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n769), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  INV_X1 U845 ( .A(G57), .ZN(G237) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U847 ( .A(n771), .B(KEYINPUT10), .ZN(n772) );
  XNOR2_X1 U848 ( .A(KEYINPUT68), .B(n772), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n837) );
  NAND2_X1 U850 ( .A1(n837), .A2(G567), .ZN(n773) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n773), .Z(G234) );
  XOR2_X1 U852 ( .A(G860), .B(KEYINPUT70), .Z(n780) );
  OR2_X1 U853 ( .A1(n780), .A2(n986), .ZN(G153) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n775) );
  INV_X1 U855 ( .A(G868), .ZN(n821) );
  NAND2_X1 U856 ( .A1(n651), .A2(n821), .ZN(n774) );
  NAND2_X1 U857 ( .A1(n775), .A2(n774), .ZN(G284) );
  NAND2_X1 U858 ( .A1(n929), .A2(n821), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT75), .ZN(n778) );
  NOR2_X1 U860 ( .A1(n821), .A2(G286), .ZN(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U862 ( .A(KEYINPUT76), .B(n779), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n781), .A2(n865), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT16), .ZN(n783) );
  XOR2_X1 U866 ( .A(KEYINPUT77), .B(n783), .Z(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n986), .ZN(n786) );
  NAND2_X1 U868 ( .A1(n865), .A2(G868), .ZN(n784) );
  NOR2_X1 U869 ( .A1(G559), .A2(n784), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G123), .A2(n520), .ZN(n787) );
  XNOR2_X1 U872 ( .A(n787), .B(KEYINPUT18), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n892), .A2(G99), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U875 ( .A1(G111), .A2(n887), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G135), .A2(n895), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n932) );
  XNOR2_X1 U879 ( .A(n932), .B(G2096), .ZN(n795) );
  INV_X1 U880 ( .A(G2100), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G80), .A2(n796), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G93), .A2(n797), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n806) );
  NAND2_X1 U885 ( .A1(G55), .A2(n800), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G67), .A2(n801), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U888 ( .A(KEYINPUT79), .B(n804), .Z(n805) );
  OR2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n820) );
  NAND2_X1 U890 ( .A1(G559), .A2(n865), .ZN(n807) );
  XOR2_X1 U891 ( .A(KEYINPUT78), .B(n807), .Z(n817) );
  XOR2_X1 U892 ( .A(n817), .B(n986), .Z(n808) );
  NOR2_X1 U893 ( .A1(G860), .A2(n808), .ZN(n809) );
  XOR2_X1 U894 ( .A(n820), .B(n809), .Z(G145) );
  XOR2_X1 U895 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n810) );
  XNOR2_X1 U896 ( .A(G305), .B(n810), .ZN(n811) );
  XNOR2_X1 U897 ( .A(G166), .B(n811), .ZN(n813) );
  XNOR2_X1 U898 ( .A(G290), .B(n929), .ZN(n812) );
  XNOR2_X1 U899 ( .A(n813), .B(n812), .ZN(n814) );
  XOR2_X1 U900 ( .A(n814), .B(n986), .Z(n815) );
  XNOR2_X1 U901 ( .A(G288), .B(n815), .ZN(n816) );
  XOR2_X1 U902 ( .A(n820), .B(n816), .Z(n864) );
  XNOR2_X1 U903 ( .A(KEYINPUT83), .B(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(n864), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G868), .ZN(n823) );
  NAND2_X1 U906 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U907 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U912 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U914 ( .A1(G120), .A2(G69), .ZN(n828) );
  XNOR2_X1 U915 ( .A(KEYINPUT84), .B(n828), .ZN(n829) );
  NOR2_X1 U916 ( .A1(G237), .A2(n829), .ZN(n830) );
  NAND2_X1 U917 ( .A1(G108), .A2(n830), .ZN(n843) );
  NAND2_X1 U918 ( .A1(n843), .A2(G567), .ZN(n835) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n831) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(n831), .Z(n832) );
  NOR2_X1 U921 ( .A1(G218), .A2(n832), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G96), .A2(n833), .ZN(n844) );
  NAND2_X1 U923 ( .A1(n844), .A2(G2106), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n835), .A2(n834), .ZN(n845) );
  NAND2_X1 U925 ( .A1(G661), .A2(G483), .ZN(n836) );
  NOR2_X1 U926 ( .A1(n845), .A2(n836), .ZN(n842) );
  NAND2_X1 U927 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n837), .ZN(G217) );
  INV_X1 U929 ( .A(G661), .ZN(n839) );
  NAND2_X1 U930 ( .A1(G2), .A2(G15), .ZN(n838) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U932 ( .A(KEYINPUT110), .B(n840), .Z(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U934 ( .A1(n842), .A2(n841), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  XNOR2_X1 U936 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  INV_X1 U942 ( .A(n845), .ZN(G319) );
  XNOR2_X1 U943 ( .A(G1986), .B(KEYINPUT41), .ZN(n855) );
  XOR2_X1 U944 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(G1981), .B(G1966), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT112), .B(G2474), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2678), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(G227) );
  XOR2_X1 U963 ( .A(n864), .B(G286), .Z(n867) );
  XNOR2_X1 U964 ( .A(G171), .B(n865), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  NOR2_X1 U966 ( .A1(G37), .A2(n868), .ZN(G397) );
  NAND2_X1 U967 ( .A1(G100), .A2(n892), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G112), .A2(n887), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G136), .A2(n895), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT114), .ZN(n875) );
  XOR2_X1 U972 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n873) );
  NAND2_X1 U973 ( .A1(G124), .A2(n520), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U977 ( .A1(n895), .A2(G142), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(KEYINPUT116), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n892), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n881), .Z(n886) );
  NAND2_X1 U982 ( .A1(G118), .A2(n887), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G130), .A2(n520), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT115), .B(n884), .Z(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n899) );
  NAND2_X1 U987 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G127), .A2(n520), .ZN(n889) );
  NAND2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n891), .B(KEYINPUT47), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G139), .A2(n895), .ZN(n896) );
  XNOR2_X1 U994 ( .A(KEYINPUT117), .B(n896), .ZN(n897) );
  NOR2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n937) );
  XOR2_X1 U996 ( .A(n899), .B(n937), .Z(n902) );
  XNOR2_X1 U997 ( .A(G164), .B(n900), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(G160), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1001 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G162), .B(n932), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(KEYINPUT118), .B(n913), .ZN(G395) );
  XOR2_X1 U1008 ( .A(KEYINPUT109), .B(G2427), .Z(n915) );
  XNOR2_X1 U1009 ( .A(G2435), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n922) );
  XOR2_X1 U1011 ( .A(G2443), .B(G2430), .Z(n917) );
  XNOR2_X1 U1012 ( .A(G2454), .B(G2446), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n918), .B(G2451), .Z(n920) );
  XNOR2_X1 U1015 ( .A(G1341), .B(G1348), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n923), .A2(G14), .ZN(n930) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n930), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n924), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G397), .A2(G395), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(n929), .ZN(G299) );
  INV_X1 U1027 ( .A(n930), .ZN(G401) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n956) );
  XOR2_X1 U1029 ( .A(G2084), .B(G160), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n950) );
  XOR2_X1 U1033 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT50), .B(n940), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT120), .ZN(n948) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(KEYINPUT51), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(n956), .B(n955), .ZN(n957) );
  OR2_X1 U1047 ( .A1(KEYINPUT55), .A2(n957), .ZN(n958) );
  NAND2_X1 U1048 ( .A1(G29), .A2(n958), .ZN(n1036) );
  XOR2_X1 U1049 ( .A(G2084), .B(KEYINPUT54), .Z(n959) );
  XNOR2_X1 U1050 ( .A(G34), .B(n959), .ZN(n976) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G35), .ZN(n974) );
  XOR2_X1 U1052 ( .A(G2072), .B(G33), .Z(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(G28), .ZN(n971) );
  XOR2_X1 U1054 ( .A(n961), .B(G27), .Z(n964) );
  XOR2_X1 U1055 ( .A(G32), .B(KEYINPUT122), .Z(n962) );
  XNOR2_X1 U1056 ( .A(n962), .B(G1996), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT123), .B(n965), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1991), .B(G25), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT53), .B(n972), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(n977), .B(KEYINPUT124), .ZN(n978) );
  XOR2_X1 U1068 ( .A(n978), .B(KEYINPUT55), .Z(n980) );
  INV_X1 U1069 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n981), .ZN(n1034) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G299), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G1341), .B(n986), .Z(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1081 ( .A(G171), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT57), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT125), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(n651), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  INV_X1 U1091 ( .A(G16), .ZN(n1030) );
  XNOR2_X1 U1092 ( .A(n1005), .B(G5), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G21), .B(G1966), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1020) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G20), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(n1017), .B(KEYINPUT60), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

