//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G155gat), .B(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n206), .A3(new_n204), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(KEYINPUT82), .A3(new_n209), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT3), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G120gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G113gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT72), .ZN(new_n217));
  INV_X1    g016(.A(G113gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n218), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT72), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n215), .B2(G113gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT71), .B1(new_n218), .B2(G120gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n218), .A2(G120gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT70), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n225), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n210), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT83), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n226), .A2(new_n232), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n234), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n234), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n237), .A2(new_n240), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT84), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n246), .B(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n212), .A2(new_n213), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n233), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT5), .A3(new_n239), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G57gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G85gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n249), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n249), .A2(KEYINPUT6), .A3(new_n261), .A4(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT24), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT65), .B1(new_n276), .B2(KEYINPUT23), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n285), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n281), .A4(new_n280), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n275), .A2(new_n288), .A3(new_n289), .A4(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n285), .A2(KEYINPUT26), .A3(new_n276), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n269), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n266), .ZN(new_n299));
  NAND2_X1  g098(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n300));
  AOI21_X1  g099(.A(G190gat), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n302));
  OAI21_X1  g101(.A(KEYINPUT68), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n300), .ZN(new_n304));
  NOR2_X1   g103(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n267), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT69), .B1(new_n304), .B2(new_n305), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n299), .A2(new_n313), .A3(new_n300), .ZN(new_n314));
  AOI211_X1 g113(.A(new_n311), .B(G190gat), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n297), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n317));
  AND2_X1   g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n317), .B1(new_n320), .B2(KEYINPUT24), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(new_n290), .A3(new_n281), .A4(new_n280), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT25), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n293), .A2(new_n316), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT69), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n299), .B2(new_n300), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT28), .B(new_n267), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(new_n303), .A3(new_n309), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(new_n297), .B1(KEYINPUT25), .B2(new_n322), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n331), .B2(new_n293), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n326), .B1(new_n332), .B2(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT77), .B(KEYINPUT22), .Z(new_n335));
  OR2_X1    g134(.A1(KEYINPUT78), .A2(G218gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT78), .A2(G218gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(G211gat), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G211gat), .A2(G218gat), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n339), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n334), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n334), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n333), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(G64gat), .ZN(new_n357));
  INV_X1    g156(.A(G92gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n333), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT81), .B1(new_n332), .B2(new_n325), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n354), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n355), .B(new_n359), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n359), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n361), .B2(new_n362), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT30), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n265), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n348), .B2(new_n349), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n250), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n348), .A2(new_n349), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n381), .A2(new_n351), .B1(new_n382), .B2(new_n236), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT86), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n346), .B2(new_n347), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n234), .B1(new_n385), .B2(new_n235), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n377), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n236), .A2(new_n382), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n352), .B2(new_n353), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n376), .A4(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT87), .ZN(new_n394));
  INV_X1    g193(.A(G22gat), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n384), .A2(new_n387), .A3(new_n395), .A4(new_n391), .ZN(new_n396));
  XNOR2_X1  g195(.A(G50gat), .B(G78gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G106gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n393), .A2(new_n394), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(KEYINPUT87), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n400), .B1(new_n393), .B2(new_n396), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n374), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT36), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n324), .A2(new_n233), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n331), .A2(new_n241), .A3(new_n293), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G227gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n410), .A2(KEYINPUT34), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n415));
  AND4_X1   g214(.A1(new_n241), .A2(new_n293), .A3(new_n316), .A4(new_n323), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n241), .B1(new_n331), .B2(new_n293), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n413), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n421), .A2(KEYINPUT75), .A3(KEYINPUT34), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT75), .B1(new_n421), .B2(KEYINPUT34), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT76), .B(new_n414), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT73), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n410), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT32), .B1(new_n429), .B2(new_n419), .ZN(new_n430));
  XOR2_X1   g229(.A(G15gat), .B(G43gat), .Z(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n419), .B1(new_n408), .B2(new_n409), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(KEYINPUT33), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n430), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n426), .A2(KEYINPUT73), .A3(new_n436), .A4(new_n427), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n407), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n426), .A2(new_n436), .A3(new_n427), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n436), .B1(new_n426), .B2(new_n427), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT36), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n406), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT88), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT37), .B(new_n355), .C1(new_n363), .C2(new_n364), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n367), .B2(new_n368), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT38), .A4(new_n359), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n361), .A2(new_n364), .A3(new_n362), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n333), .A2(new_n354), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT37), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT90), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT37), .A4(new_n451), .ZN(new_n455));
  AND4_X1   g254(.A1(new_n359), .A2(new_n453), .A3(new_n448), .A4(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n449), .B1(new_n456), .B2(KEYINPUT38), .ZN(new_n457));
  INV_X1    g256(.A(new_n265), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n369), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n403), .A2(new_n400), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n393), .A2(new_n396), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n401), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  INV_X1    g263(.A(new_n237), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n244), .A2(new_n245), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n239), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n261), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n467), .B(KEYINPUT39), .C1(new_n239), .C2(new_n252), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(KEYINPUT89), .A3(KEYINPUT40), .A4(new_n470), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n373), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n472), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n262), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n463), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n406), .C1(new_n440), .C2(new_n443), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n445), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n424), .A2(new_n425), .ZN(new_n483));
  INV_X1    g282(.A(new_n427), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n437), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n426), .A2(new_n436), .A3(new_n427), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n405), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  INV_X1    g287(.A(new_n374), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n487), .A2(KEYINPUT91), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n488), .B(new_n463), .C1(new_n441), .C2(new_n442), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n374), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n405), .B(new_n374), .C1(new_n439), .C2(new_n438), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n490), .B(new_n493), .C1(new_n494), .C2(new_n488), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n482), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT14), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G43gat), .ZN(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(KEYINPUT93), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT93), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n497), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n504), .B2(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT93), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n522), .A2(new_n523), .B1(new_n511), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n532), .B2(KEYINPUT94), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(G1gat), .B2(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI221_X1 g334(.A(new_n532), .B1(KEYINPUT94), .B2(new_n528), .C1(G1gat), .C2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n519), .B2(new_n518), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n518), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n537), .B(new_n525), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n541), .B(KEYINPUT13), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n527), .A2(new_n538), .B1(new_n537), .B2(new_n518), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n541), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G169gat), .B(G197gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT96), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n550), .A2(KEYINPUT96), .A3(new_n557), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n544), .A2(new_n547), .A3(new_n549), .A4(new_n556), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  OAI22_X1  g362(.A1(new_n558), .A2(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G190gat), .B(G218gat), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n518), .A2(new_n519), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n358), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n569), .B2(new_n358), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n575), .A3(new_n572), .A4(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT100), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n527), .A2(new_n567), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585));
  AND2_X1   g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n582), .A2(new_n518), .B1(KEYINPUT41), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n566), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI221_X4 g389(.A(new_n582), .B1(new_n519), .B2(new_n518), .C1(new_n520), .C2(new_n526), .ZN(new_n591));
  INV_X1    g390(.A(new_n587), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT101), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n565), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n586), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n596), .B1(new_n590), .B2(new_n595), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  OR2_X1    g404(.A1(G57gat), .A2(G64gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(G57gat), .A2(G64gat), .ZN(new_n607));
  AND2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(KEYINPUT9), .ZN(new_n609));
  NOR2_X1   g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(KEYINPUT98), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n608), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n609), .B(new_n611), .C1(new_n608), .C2(new_n610), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n614), .A2(new_n615), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n537), .B1(KEYINPUT21), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n266), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n616), .A2(new_n617), .ZN(new_n626));
  OAI21_X1  g425(.A(G183gat), .B1(new_n626), .B2(new_n537), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n627), .A3(new_n622), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n629), .A2(G231gat), .A3(G233gat), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n628), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n340), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n631), .B2(new_n634), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n621), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n620), .A3(new_n638), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n614), .A2(new_n615), .B1(new_n577), .B2(new_n578), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n582), .B2(new_n616), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n284), .ZN(new_n651));
  INV_X1    g450(.A(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n582), .A2(KEYINPUT10), .A3(new_n623), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n646), .B2(KEYINPUT10), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n656), .A2(KEYINPUT103), .A3(new_n647), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT103), .B1(new_n656), .B2(new_n647), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n649), .B(new_n654), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n647), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n649), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n653), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n605), .A2(new_n644), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT104), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667));
  NOR4_X1   g466(.A1(new_n605), .A2(new_n644), .A3(new_n667), .A4(new_n664), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n496), .A2(new_n564), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n458), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g471(.A(new_n528), .B1(new_n670), .B2(new_n476), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n496), .A2(new_n564), .A3(new_n669), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(G8gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n530), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n674), .A2(new_n373), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n679), .B(new_n680), .C1(KEYINPUT42), .C2(new_n678), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n670), .A2(new_n476), .A3(new_n676), .ZN(new_n683));
  OAI21_X1  g482(.A(G8gat), .B1(new_n674), .B2(new_n373), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT106), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(G1325gat));
  NOR2_X1   g487(.A1(new_n441), .A2(new_n442), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(G15gat), .B1(new_n670), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n440), .A2(new_n443), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT107), .B1(new_n440), .B2(new_n443), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n674), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n691), .B1(G15gat), .B2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n674), .A2(new_n463), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n590), .A2(new_n595), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n597), .A3(new_n600), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n597), .B2(new_n600), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n479), .B(new_n406), .C1(new_n440), .C2(new_n443), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n495), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n482), .B2(new_n495), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n644), .ZN(new_n714));
  INV_X1    g513(.A(new_n558), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n550), .A2(KEYINPUT96), .A3(new_n557), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n542), .A2(new_n543), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT18), .B1(new_n548), .B2(new_n541), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(KEYINPUT97), .A3(new_n547), .A4(new_n556), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n560), .A2(new_n561), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n715), .A2(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n714), .A2(new_n722), .A3(new_n664), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n713), .A2(new_n458), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n711), .A2(new_n498), .A3(new_n458), .A4(new_n723), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT110), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(G29gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n729), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(G1328gat));
  NAND2_X1  g534(.A1(new_n711), .A2(new_n723), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(G36gat), .A3(new_n373), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n713), .A2(new_n476), .A3(new_n723), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n499), .B2(new_n739), .ZN(G1329gat));
  NAND4_X1  g539(.A1(new_n711), .A2(new_n507), .A3(new_n690), .A4(new_n723), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n713), .A2(new_n692), .A3(new_n723), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT47), .B(new_n741), .C1(new_n742), .C2(new_n507), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n713), .A2(new_n696), .A3(new_n723), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n741), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g546(.A(new_n505), .B1(new_n736), .B2(new_n463), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n713), .A2(G50gat), .A3(new_n723), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n463), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT48), .ZN(G1331gat));
  AOI211_X1 g550(.A(new_n644), .B(new_n605), .C1(new_n495), .C2(new_n707), .ZN(new_n752));
  INV_X1    g551(.A(new_n664), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n564), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n458), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g556(.A1(new_n752), .A2(new_n754), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n373), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n758), .B2(new_n697), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(new_n690), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(G71gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n758), .A2(new_n463), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(G78gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT112), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n769), .B(new_n771), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n714), .A2(new_n564), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n708), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT113), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n265), .A2(G85gat), .A3(new_n753), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n773), .A2(new_n664), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n713), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n458), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G85gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n790), .ZN(G1336gat));
  AOI21_X1  g590(.A(new_n712), .B1(new_n496), .B2(new_n605), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n495), .A2(new_n707), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(new_n605), .A3(new_n709), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n476), .B(new_n787), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n373), .A2(G92gat), .A3(new_n753), .ZN(new_n797));
  AND4_X1   g596(.A1(KEYINPUT51), .A2(new_n793), .A3(new_n605), .A4(new_n773), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n708), .B2(new_n773), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n796), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  INV_X1    g605(.A(new_n797), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n796), .B(new_n806), .C1(new_n780), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1337gat));
  NOR3_X1   g608(.A1(new_n689), .A2(G99gat), .A3(new_n753), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n781), .A2(new_n783), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n788), .A2(new_n696), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G99gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1338gat));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n463), .A2(G106gat), .A3(new_n753), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n780), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n713), .A2(new_n405), .A3(new_n787), .ZN(new_n818));
  XOR2_X1   g617(.A(KEYINPUT116), .B(G106gat), .Z(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n816), .B1(new_n776), .B2(new_n777), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n818), .B2(new_n820), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n817), .A2(new_n821), .B1(new_n823), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g623(.A(new_n659), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n653), .B1(new_n660), .B2(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n648), .B(new_n655), .C1(new_n646), .C2(KEYINPUT10), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n827), .B2(KEYINPUT117), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT103), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n660), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n656), .A2(KEYINPUT103), .A3(new_n647), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n825), .B1(new_n834), .B2(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n834), .B2(KEYINPUT55), .ZN(new_n837));
  INV_X1    g636(.A(new_n826), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n646), .A2(KEYINPUT10), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n648), .A4(new_n655), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT54), .B(new_n841), .C1(new_n657), .C2(new_n658), .ZN(new_n842));
  INV_X1    g641(.A(new_n833), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n564), .A2(new_n835), .A3(new_n837), .A4(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n555), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n548), .A2(new_n541), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n545), .A2(new_n546), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n720), .B2(new_n721), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n664), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n605), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n852), .A2(new_n837), .A3(new_n835), .A4(new_n846), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n706), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n644), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n665), .A2(new_n722), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n476), .A2(new_n265), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n438), .A2(new_n439), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n463), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n218), .A3(new_n564), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n859), .A2(new_n487), .A3(new_n860), .ZN(new_n866));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n722), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1340gat));
  OAI21_X1  g667(.A(G120gat), .B1(new_n866), .B2(new_n753), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT119), .Z(new_n870));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n215), .A3(new_n664), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n866), .A2(new_n873), .A3(new_n644), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n864), .A2(new_n714), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n873), .ZN(G1342gat));
  INV_X1    g675(.A(G134gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n864), .A2(new_n877), .A3(new_n605), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT56), .Z(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n866), .B2(new_n706), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n861), .A2(new_n696), .A3(new_n463), .ZN(new_n886));
  INV_X1    g685(.A(G141gat), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n564), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n844), .A2(new_n845), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT55), .B(new_n838), .C1(new_n842), .C2(new_n843), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n659), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n853), .B1(new_n722), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n706), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n837), .A2(new_n846), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n605), .A2(new_n895), .A3(new_n835), .A4(new_n852), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n714), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n858), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n559), .A2(new_n558), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n560), .B(KEYINPUT97), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n835), .B(new_n890), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n605), .B1(new_n901), .B2(new_n853), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT121), .B(new_n644), .C1(new_n902), .C2(new_n856), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n405), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n860), .B1(new_n440), .B2(new_n443), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n463), .B1(new_n857), .B2(new_n858), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n889), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n644), .B1(new_n902), .B2(new_n856), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n858), .A3(new_n903), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n909), .B1(new_n915), .B2(new_n405), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n837), .A2(new_n835), .A3(new_n846), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n853), .B1(new_n917), .B2(new_n722), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n706), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n714), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n665), .A2(new_n722), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n909), .B(new_n405), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n907), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n916), .A2(KEYINPUT122), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n564), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n888), .B1(new_n926), .B2(G141gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n916), .A2(new_n924), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n887), .B1(new_n929), .B2(new_n564), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n927), .A2(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1344gat));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n859), .A2(new_n405), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT57), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n666), .A2(new_n668), .A3(new_n564), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n909), .B(new_n405), .C1(new_n936), .C2(new_n897), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n937), .A3(new_n664), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n933), .B1(new_n938), .B2(new_n907), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G148gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n938), .A2(new_n933), .A3(new_n907), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT59), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n664), .B1(new_n911), .B2(new_n925), .ZN(new_n944));
  INV_X1    g743(.A(G148gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT59), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT122), .B1(new_n916), .B2(new_n924), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n921), .B1(new_n912), .B2(new_n913), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n463), .B1(new_n949), .B2(new_n903), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n910), .B(new_n889), .C1(new_n950), .C2(new_n909), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n753), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n946), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(KEYINPUT123), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n942), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n886), .A2(new_n945), .A3(new_n664), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1345gat));
  AOI21_X1  g756(.A(G155gat), .B1(new_n886), .B2(new_n714), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n644), .B1(new_n948), .B2(new_n951), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g759(.A(G162gat), .B1(new_n886), .B2(new_n605), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n706), .B1(new_n948), .B2(new_n951), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(G162gat), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n458), .B1(new_n857), .B2(new_n858), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n476), .A3(new_n487), .ZN(new_n965));
  OAI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n722), .ZN(new_n966));
  AOI211_X1 g765(.A(new_n458), .B(new_n863), .C1(new_n857), .C2(new_n858), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n476), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n564), .A2(new_n283), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1348gat));
  NOR3_X1   g769(.A1(new_n965), .A2(new_n284), .A3(new_n753), .ZN(new_n971));
  INV_X1    g770(.A(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n664), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n973), .B2(new_n284), .ZN(G1349gat));
  NOR2_X1   g773(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n972), .B(new_n714), .C1(new_n328), .C2(new_n327), .ZN(new_n976));
  OAI21_X1  g775(.A(G183gat), .B1(new_n965), .B2(new_n644), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n978), .B(new_n979), .Z(G1350gat));
  NAND3_X1  g779(.A1(new_n972), .A2(new_n267), .A3(new_n605), .ZN(new_n981));
  OAI21_X1  g780(.A(G190gat), .B1(new_n965), .B2(new_n706), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1351gat));
  NOR2_X1   g784(.A1(new_n696), .A2(new_n373), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(new_n405), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n989), .A3(new_n405), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n988), .A2(new_n964), .A3(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(G197gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n992), .A2(new_n993), .A3(new_n564), .ZN(new_n994));
  AND4_X1   g793(.A1(new_n265), .A2(new_n986), .A3(new_n935), .A4(new_n937), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n995), .A2(new_n564), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n994), .B1(new_n993), .B2(new_n996), .ZN(G1352gat));
  NAND3_X1  g796(.A1(new_n992), .A2(new_n652), .A3(new_n664), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n986), .A2(new_n265), .ZN(new_n1000));
  OAI21_X1  g799(.A(G204gat), .B1(new_n938), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n992), .A2(new_n1002), .A3(new_n652), .A4(new_n664), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(G1353gat));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n991), .A2(new_n644), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1005), .B1(new_n1006), .B2(new_n340), .ZN(new_n1007));
  NOR4_X1   g806(.A1(new_n991), .A2(KEYINPUT127), .A3(G211gat), .A4(new_n644), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n995), .A2(new_n714), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1009), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT63), .B1(new_n1009), .B2(G211gat), .ZN(new_n1011));
  OAI22_X1  g810(.A1(new_n1007), .A2(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  AND4_X1   g811(.A1(new_n605), .A2(new_n995), .A3(new_n336), .A4(new_n337), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n992), .A2(new_n605), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1013), .B1(new_n1014), .B2(new_n341), .ZN(G1355gat));
endmodule


