

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U557 ( .A1(G160), .A2(n597), .ZN(n664) );
  BUF_X1 U558 ( .A(n712), .Z(n713) );
  NOR2_X1 U559 ( .A1(n577), .A2(G651), .ZN(n525) );
  NOR2_X1 U560 ( .A1(n551), .A2(G2104), .ZN(n546) );
  XNOR2_X1 U561 ( .A(n545), .B(n544), .ZN(n548) );
  XNOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n544) );
  NOR2_X1 U563 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n788) );
  INV_X1 U565 ( .A(KEYINPUT68), .ZN(n549) );
  XOR2_X2 U566 ( .A(KEYINPUT65), .B(n525), .Z(n526) );
  INV_X1 U567 ( .A(G2105), .ZN(n551) );
  NAND2_X1 U568 ( .A1(G160), .A2(G40), .ZN(n523) );
  XOR2_X1 U569 ( .A(n646), .B(KEYINPUT28), .Z(n524) );
  INV_X1 U570 ( .A(KEYINPUT91), .ZN(n624) );
  XNOR2_X1 U571 ( .A(n625), .B(n624), .ZN(n626) );
  INV_X1 U572 ( .A(KEYINPUT29), .ZN(n648) );
  INV_X1 U573 ( .A(KEYINPUT31), .ZN(n660) );
  XNOR2_X1 U574 ( .A(n661), .B(n660), .ZN(n662) );
  INV_X1 U575 ( .A(n921), .ZN(n692) );
  NOR2_X1 U576 ( .A1(n693), .A2(n692), .ZN(n694) );
  INV_X1 U577 ( .A(G651), .ZN(n535) );
  INV_X1 U578 ( .A(G2105), .ZN(n543) );
  NOR2_X1 U579 ( .A1(n711), .A2(n710), .ZN(n745) );
  AND2_X1 U580 ( .A1(n543), .A2(G2104), .ZN(n883) );
  XNOR2_X1 U581 ( .A(KEYINPUT70), .B(n529), .ZN(n785) );
  XNOR2_X1 U582 ( .A(KEYINPUT76), .B(n542), .ZN(G168) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NAND2_X1 U584 ( .A1(n526), .A2(G51), .ZN(n527) );
  XOR2_X1 U585 ( .A(KEYINPUT75), .B(n527), .Z(n531) );
  NOR2_X1 U586 ( .A1(G543), .A2(n535), .ZN(n528) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n528), .Z(n529) );
  NAND2_X1 U588 ( .A1(G63), .A2(n785), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U590 ( .A(KEYINPUT6), .B(n532), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G89), .A2(n788), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n533), .B(KEYINPUT4), .ZN(n534) );
  XNOR2_X1 U593 ( .A(n534), .B(KEYINPUT74), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n577), .A2(n535), .ZN(n789) );
  NAND2_X1 U595 ( .A1(G76), .A2(n789), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U597 ( .A(n538), .B(KEYINPUT5), .Z(n539) );
  NOR2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U599 ( .A(n541), .B(KEYINPUT7), .Z(n542) );
  NAND2_X1 U600 ( .A1(G101), .A2(n883), .ZN(n545) );
  XNOR2_X2 U601 ( .A(n546), .B(KEYINPUT66), .ZN(n886) );
  NAND2_X1 U602 ( .A1(G125), .A2(n886), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U604 ( .A(n550), .B(n549), .ZN(n553) );
  AND2_X1 U605 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U606 ( .A1(n888), .A2(G113), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n557) );
  NOR2_X1 U608 ( .A1(G2105), .A2(G2104), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT17), .B(n554), .Z(n712) );
  NAND2_X1 U610 ( .A1(G137), .A2(n712), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT69), .B(n555), .ZN(n556) );
  NOR2_X2 U612 ( .A1(n557), .A2(n556), .ZN(G160) );
  NAND2_X1 U613 ( .A1(G102), .A2(n883), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G138), .A2(n712), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G114), .A2(n888), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G126), .A2(n886), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(G164) );
  NAND2_X1 U620 ( .A1(n526), .A2(G52), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G64), .A2(n785), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G90), .A2(n788), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G77), .A2(n789), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U627 ( .A1(n570), .A2(n569), .ZN(G171) );
  XOR2_X1 U628 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U629 ( .A1(G88), .A2(n788), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G75), .A2(n789), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n526), .A2(G50), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G62), .A2(n785), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U635 ( .A1(n576), .A2(n575), .ZN(G166) );
  INV_X1 U636 ( .A(G166), .ZN(G303) );
  NAND2_X1 U637 ( .A1(G49), .A2(n526), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n785), .A2(n580), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G651), .A2(G74), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G73), .A2(n789), .ZN(n583) );
  XNOR2_X1 U644 ( .A(n583), .B(KEYINPUT2), .ZN(n590) );
  NAND2_X1 U645 ( .A1(G86), .A2(n788), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G61), .A2(n785), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G48), .A2(n526), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT79), .B(n586), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G85), .A2(n788), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G72), .A2(n789), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U655 ( .A1(n526), .A2(G47), .ZN(n594) );
  NAND2_X1 U656 ( .A1(G60), .A2(n785), .ZN(n593) );
  NAND2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U658 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n709) );
  AND2_X1 U660 ( .A1(n709), .A2(G40), .ZN(n597) );
  AND2_X1 U661 ( .A1(n664), .A2(G1341), .ZN(n609) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n788), .A2(G81), .ZN(n598) );
  XNOR2_X1 U664 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G68), .A2(n789), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n602), .B(n601), .ZN(n606) );
  NAND2_X1 U668 ( .A1(G56), .A2(n785), .ZN(n603) );
  XNOR2_X1 U669 ( .A(KEYINPUT14), .B(n603), .ZN(n604) );
  INV_X1 U670 ( .A(n604), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U672 ( .A1(n526), .A2(G43), .ZN(n607) );
  NAND2_X1 U673 ( .A1(n608), .A2(n607), .ZN(n933) );
  NOR2_X1 U674 ( .A1(n609), .A2(n933), .ZN(n613) );
  XNOR2_X1 U675 ( .A(G1996), .B(KEYINPUT89), .ZN(n944) );
  NOR2_X1 U676 ( .A1(n664), .A2(n944), .ZN(n611) );
  XOR2_X1 U677 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n612) );
  AND2_X1 U679 ( .A1(n613), .A2(n612), .ZN(n631) );
  NAND2_X1 U680 ( .A1(G54), .A2(n526), .ZN(n620) );
  NAND2_X1 U681 ( .A1(G79), .A2(n789), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G66), .A2(n785), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G92), .A2(n788), .ZN(n616) );
  XNOR2_X1 U685 ( .A(KEYINPUT73), .B(n616), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n621), .B(KEYINPUT15), .ZN(n924) );
  NAND2_X1 U689 ( .A1(n631), .A2(n924), .ZN(n630) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n664), .ZN(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT90), .B(n622), .ZN(n627) );
  INV_X1 U692 ( .A(n664), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n623), .A2(G2067), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT92), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n633) );
  OR2_X1 U697 ( .A1(n924), .A2(n631), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n644) );
  NAND2_X1 U699 ( .A1(n623), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  AND2_X1 U701 ( .A1(G1956), .A2(n664), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n645) );
  NAND2_X1 U703 ( .A1(n526), .A2(G53), .ZN(n638) );
  NAND2_X1 U704 ( .A1(G65), .A2(n785), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U706 ( .A1(G91), .A2(n788), .ZN(n640) );
  NAND2_X1 U707 ( .A1(G78), .A2(n789), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n934) );
  NAND2_X1 U710 ( .A1(n645), .A2(n934), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n645), .A2(n934), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n647), .A2(n524), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n653) );
  INV_X1 U715 ( .A(G1961), .ZN(n971) );
  NAND2_X1 U716 ( .A1(n664), .A2(n971), .ZN(n651) );
  XNOR2_X1 U717 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U718 ( .A1(n623), .A2(n945), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U720 ( .A1(n657), .A2(G171), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n663) );
  NAND2_X1 U722 ( .A1(G8), .A2(n664), .ZN(n704) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n704), .ZN(n677) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n664), .ZN(n674) );
  NOR2_X1 U725 ( .A1(n677), .A2(n674), .ZN(n654) );
  NAND2_X1 U726 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U728 ( .A1(G168), .A2(n656), .ZN(n659) );
  NOR2_X1 U729 ( .A1(G171), .A2(n657), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n675) );
  NAND2_X1 U731 ( .A1(n675), .A2(G286), .ZN(n670) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n704), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT93), .B(n667), .Z(n668) );
  NAND2_X1 U736 ( .A1(n668), .A2(G303), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n671), .B(KEYINPUT94), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n672), .A2(G8), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT32), .ZN(n681) );
  NAND2_X1 U741 ( .A1(G8), .A2(n674), .ZN(n679) );
  INV_X1 U742 ( .A(n675), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n699) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n918) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n918), .A2(n682), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n699), .A2(n683), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT95), .ZN(n688) );
  NAND2_X1 U751 ( .A1(G288), .A2(G1976), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n685), .B(KEYINPUT96), .ZN(n925) );
  INV_X1 U753 ( .A(n925), .ZN(n686) );
  OR2_X1 U754 ( .A1(n686), .A2(n704), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n689), .A2(KEYINPUT33), .ZN(n690) );
  INV_X1 U757 ( .A(n690), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n918), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n691), .A2(n704), .ZN(n693) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT97), .ZN(n708) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U764 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n704), .A2(n700), .ZN(n706) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n701) );
  XOR2_X1 U768 ( .A(n701), .B(KEYINPUT88), .Z(n702) );
  XNOR2_X1 U769 ( .A(KEYINPUT24), .B(n702), .ZN(n703) );
  OR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n711) );
  XNOR2_X1 U773 ( .A(G1986), .B(G290), .ZN(n938) );
  NOR2_X1 U774 ( .A1(n709), .A2(n523), .ZN(n756) );
  AND2_X1 U775 ( .A1(n938), .A2(n756), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n724) );
  NAND2_X1 U777 ( .A1(G104), .A2(n883), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G140), .A2(n713), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U780 ( .A(KEYINPUT34), .B(n716), .ZN(n721) );
  NAND2_X1 U781 ( .A1(G116), .A2(n888), .ZN(n718) );
  NAND2_X1 U782 ( .A1(G128), .A2(n886), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U784 ( .A(n719), .B(KEYINPUT35), .Z(n720) );
  NOR2_X1 U785 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U786 ( .A(KEYINPUT84), .B(n722), .Z(n723) );
  XNOR2_X1 U787 ( .A(n724), .B(n723), .ZN(n899) );
  XNOR2_X1 U788 ( .A(KEYINPUT37), .B(G2067), .ZN(n754) );
  NOR2_X1 U789 ( .A1(n899), .A2(n754), .ZN(n725) );
  XNOR2_X1 U790 ( .A(KEYINPUT86), .B(n725), .ZN(n1005) );
  NAND2_X1 U791 ( .A1(n756), .A2(n1005), .ZN(n752) );
  NAND2_X1 U792 ( .A1(G117), .A2(n888), .ZN(n727) );
  NAND2_X1 U793 ( .A1(G129), .A2(n886), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U795 ( .A1(n883), .A2(G105), .ZN(n728) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n728), .Z(n729) );
  NOR2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U798 ( .A1(n713), .A2(G141), .ZN(n731) );
  NAND2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n868) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n868), .ZN(n733) );
  XNOR2_X1 U801 ( .A(n733), .B(KEYINPUT87), .ZN(n741) );
  INV_X1 U802 ( .A(G1991), .ZN(n746) );
  NAND2_X1 U803 ( .A1(G95), .A2(n883), .ZN(n735) );
  NAND2_X1 U804 ( .A1(G107), .A2(n888), .ZN(n734) );
  NAND2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U806 ( .A1(G131), .A2(n713), .ZN(n737) );
  NAND2_X1 U807 ( .A1(G119), .A2(n886), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n898) );
  NOR2_X1 U810 ( .A1(n746), .A2(n898), .ZN(n740) );
  NOR2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n1013) );
  INV_X1 U812 ( .A(n756), .ZN(n742) );
  NOR2_X1 U813 ( .A1(n1013), .A2(n742), .ZN(n749) );
  INV_X1 U814 ( .A(n749), .ZN(n743) );
  AND2_X1 U815 ( .A1(n752), .A2(n743), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n759) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n868), .ZN(n1010) );
  AND2_X1 U818 ( .A1(n746), .A2(n898), .ZN(n1003) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U820 ( .A1(n1003), .A2(n747), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U822 ( .A1(n1010), .A2(n750), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U825 ( .A1(n899), .A2(n754), .ZN(n1012) );
  NAND2_X1 U826 ( .A1(n755), .A2(n1012), .ZN(n757) );
  NAND2_X1 U827 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U829 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U831 ( .A(G132), .ZN(G219) );
  INV_X1 U832 ( .A(G82), .ZN(G220) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n821) );
  NAND2_X1 U837 ( .A1(n821), .A2(G567), .ZN(n762) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  XOR2_X1 U839 ( .A(G860), .B(KEYINPUT72), .Z(n768) );
  OR2_X1 U840 ( .A1(n768), .A2(n933), .ZN(G153) );
  INV_X1 U841 ( .A(G171), .ZN(G301) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n764) );
  OR2_X1 U843 ( .A1(n924), .A2(G868), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n764), .A2(n763), .ZN(G284) );
  INV_X1 U845 ( .A(n934), .ZN(G299) );
  XNOR2_X1 U846 ( .A(KEYINPUT77), .B(G868), .ZN(n765) );
  NOR2_X1 U847 ( .A1(G286), .A2(n765), .ZN(n767) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U849 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n768), .A2(G559), .ZN(n769) );
  NAND2_X1 U851 ( .A1(n769), .A2(n924), .ZN(n770) );
  XNOR2_X1 U852 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G868), .A2(n933), .ZN(n773) );
  NAND2_X1 U854 ( .A1(G868), .A2(n924), .ZN(n771) );
  NOR2_X1 U855 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U856 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U857 ( .A1(G99), .A2(n883), .ZN(n775) );
  NAND2_X1 U858 ( .A1(G111), .A2(n888), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n780) );
  NAND2_X1 U860 ( .A1(n886), .A2(G123), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT18), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n713), .A2(G135), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n1004) );
  XNOR2_X1 U865 ( .A(n1004), .B(G2096), .ZN(n781) );
  XNOR2_X1 U866 ( .A(n781), .B(KEYINPUT78), .ZN(n783) );
  INV_X1 U867 ( .A(G2100), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U869 ( .A1(G559), .A2(n924), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(n933), .ZN(n802) );
  NOR2_X1 U871 ( .A1(n802), .A2(G860), .ZN(n794) );
  NAND2_X1 U872 ( .A1(n526), .A2(G55), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G67), .A2(n785), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U875 ( .A1(G93), .A2(n788), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G80), .A2(n789), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n796) );
  XNOR2_X1 U879 ( .A(n794), .B(n796), .ZN(G145) );
  NOR2_X1 U880 ( .A1(n796), .A2(G868), .ZN(n795) );
  XNOR2_X1 U881 ( .A(KEYINPUT81), .B(n795), .ZN(n806) );
  XNOR2_X1 U882 ( .A(G166), .B(G290), .ZN(n799) );
  XNOR2_X1 U883 ( .A(n934), .B(n796), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(G305), .ZN(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U886 ( .A(KEYINPUT19), .B(n800), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(G288), .ZN(n906) );
  XNOR2_X1 U888 ( .A(n906), .B(n802), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n803), .A2(G868), .ZN(n804) );
  XNOR2_X1 U890 ( .A(KEYINPUT80), .B(n804), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n807) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n807), .Z(n808) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n808), .ZN(n809) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n809), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n810), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U898 ( .A1(G69), .A2(G120), .ZN(n811) );
  NOR2_X1 U899 ( .A1(G237), .A2(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G108), .A2(n812), .ZN(n825) );
  NAND2_X1 U901 ( .A1(n825), .A2(G567), .ZN(n818) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n813) );
  XNOR2_X1 U903 ( .A(KEYINPUT22), .B(n813), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(G96), .ZN(n815) );
  NOR2_X1 U905 ( .A1(G218), .A2(n815), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT82), .B(n816), .Z(n826) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n826), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n838) );
  NAND2_X1 U909 ( .A1(G661), .A2(G483), .ZN(n819) );
  XOR2_X1 U910 ( .A(KEYINPUT83), .B(n819), .Z(n820) );
  NOR2_X1 U911 ( .A1(n838), .A2(n820), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U924 ( .A(G2454), .B(G2451), .ZN(n835) );
  XNOR2_X1 U925 ( .A(G2430), .B(G2446), .ZN(n833) );
  XOR2_X1 U926 ( .A(G2435), .B(G2427), .Z(n828) );
  XNOR2_X1 U927 ( .A(KEYINPUT98), .B(G2438), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U929 ( .A(n829), .B(G2443), .Z(n831) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U934 ( .A1(n836), .A2(G14), .ZN(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT99), .B(n837), .ZN(n915) );
  XNOR2_X1 U936 ( .A(n915), .B(KEYINPUT100), .ZN(G401) );
  INV_X1 U937 ( .A(n838), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2090), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2072), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n841), .B(G2096), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2084), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2678), .Z(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT101), .B(G2100), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G1976), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1961), .B(G1956), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n850), .B(KEYINPUT103), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(G1981), .B(G1971), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT102), .B(G2474), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G100), .A2(n883), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G112), .A2(n888), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n867) );
  NAND2_X1 U963 ( .A1(n886), .A2(G124), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n861), .B(KEYINPUT104), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G136), .A2(n713), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT105), .B(n865), .Z(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U970 ( .A(n868), .B(G162), .ZN(n870) );
  XNOR2_X1 U971 ( .A(G164), .B(G160), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n882) );
  NAND2_X1 U973 ( .A1(n886), .A2(G130), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(KEYINPUT106), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G118), .A2(n888), .ZN(n872) );
  XOR2_X1 U976 ( .A(KEYINPUT107), .B(n872), .Z(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n713), .A2(G142), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n875), .B(KEYINPUT108), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G106), .A2(n883), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(n882), .B(n881), .Z(n904) );
  NAND2_X1 U985 ( .A1(G103), .A2(n883), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G139), .A2(n713), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G127), .A2(n886), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n887), .B(KEYINPUT110), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G115), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n894), .Z(n1014) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(n897), .B(n1004), .Z(n901) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n1014), .B(n902), .Z(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n924), .B(G286), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n933), .B(G171), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G397) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(G16), .B(KEYINPUT56), .ZN(n942) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT121), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G168), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT57), .B(n923), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n924), .B(G1348), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G1971), .B(G303), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n940) );
  XOR2_X1 U1031 ( .A(n933), .B(G1341), .Z(n936) );
  XNOR2_X1 U1032 ( .A(n934), .B(G1956), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT122), .B(n943), .ZN(n1000) );
  XNOR2_X1 U1038 ( .A(n944), .B(G32), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n945), .B(G27), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT119), .B(n948), .ZN(n958) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(KEYINPUT116), .ZN(n952) );
  XOR2_X1 U1044 ( .A(G2072), .B(G33), .Z(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT117), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(KEYINPUT118), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(G28), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G25), .B(G1991), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1056 ( .A(KEYINPUT115), .B(G2090), .Z(n963) );
  XNOR2_X1 U1057 ( .A(G35), .B(n963), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n966), .ZN(n968) );
  INV_X1 U1060 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(G11), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n970), .B(KEYINPUT120), .ZN(n998) );
  XNOR2_X1 U1064 ( .A(n971), .B(G5), .ZN(n993) );
  XOR2_X1 U1065 ( .A(G1966), .B(G21), .Z(n984) );
  XNOR2_X1 U1066 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n972), .B(G4), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n973), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G6), .B(G1981), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT123), .B(n976), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT125), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n982), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n994), .B(KEYINPUT61), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT126), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n996), .A2(G16), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT127), .ZN(n1029) );
  XOR2_X1 U1093 ( .A(G160), .B(G2084), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT114), .B(n1008), .ZN(n1023) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1011), .Z(n1021) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1014), .Z(n1016) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1017), .Z(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  INV_X1 U1110 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

