

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782;

  NAND2_X1 U366 ( .A1(n576), .A2(n550), .ZN(n707) );
  XNOR2_X1 U367 ( .A(n600), .B(KEYINPUT1), .ZN(n714) );
  XOR2_X1 U368 ( .A(G122), .B(G104), .Z(n370) );
  XNOR2_X1 U369 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n492) );
  BUF_X1 U370 ( .A(n641), .Z(n694) );
  XNOR2_X2 U371 ( .A(n412), .B(KEYINPUT41), .ZN(n734) );
  NAND2_X2 U372 ( .A1(n528), .A2(G214), .ZN(n704) );
  XNOR2_X2 U373 ( .A(n650), .B(KEYINPUT93), .ZN(n751) );
  OR2_X1 U374 ( .A1(n687), .A2(n592), .ZN(n577) );
  XNOR2_X1 U375 ( .A(G143), .B(G113), .ZN(n497) );
  NOR2_X1 U376 ( .A1(n656), .A2(G902), .ZN(n505) );
  XOR2_X1 U377 ( .A(n415), .B(n467), .Z(n345) );
  XOR2_X1 U378 ( .A(n408), .B(KEYINPUT30), .Z(n346) );
  NOR2_X2 U379 ( .A1(n576), .A2(n575), .ZN(n592) );
  NAND2_X1 U380 ( .A1(n636), .A2(n635), .ZN(n769) );
  NOR2_X1 U381 ( .A1(n626), .A2(n403), .ZN(n690) );
  NAND2_X1 U382 ( .A1(n446), .A2(n443), .ZN(n711) );
  AND2_X1 U383 ( .A1(n400), .A2(n622), .ZN(n627) );
  AND2_X2 U384 ( .A1(n612), .A2(n611), .ZN(n613) );
  AND2_X1 U385 ( .A1(n374), .A2(n346), .ZN(n390) );
  XNOR2_X1 U386 ( .A(n423), .B(KEYINPUT28), .ZN(n612) );
  NOR2_X1 U387 ( .A1(n618), .A2(n719), .ZN(n423) );
  XNOR2_X1 U388 ( .A(n348), .B(KEYINPUT19), .ZN(n609) );
  NAND2_X1 U389 ( .A1(n705), .A2(n704), .ZN(n701) );
  OR2_X1 U390 ( .A1(n713), .A2(n535), .ZN(n447) );
  NAND2_X1 U391 ( .A1(n538), .A2(n704), .ZN(n348) );
  AND2_X1 U392 ( .A1(n365), .A2(n361), .ZN(n360) );
  BUF_X1 U393 ( .A(n534), .Z(n719) );
  XNOR2_X1 U394 ( .A(n413), .B(n383), .ZN(n748) );
  NAND2_X1 U395 ( .A1(n364), .A2(KEYINPUT60), .ZN(n356) );
  OR2_X1 U396 ( .A1(n364), .A2(KEYINPUT60), .ZN(n353) );
  INV_X1 U397 ( .A(n751), .ZN(n364) );
  XNOR2_X1 U398 ( .A(n507), .B(n470), .ZN(n766) );
  XOR2_X1 U399 ( .A(G131), .B(G140), .Z(n501) );
  XOR2_X1 U400 ( .A(KEYINPUT82), .B(KEYINPUT34), .Z(n458) );
  NOR2_X2 U401 ( .A1(n651), .A2(n751), .ZN(n652) );
  XNOR2_X2 U402 ( .A(n347), .B(n544), .ZN(n554) );
  NAND2_X1 U403 ( .A1(n609), .A2(n543), .ZN(n347) );
  NOR2_X1 U404 ( .A1(n742), .A2(n657), .ZN(n362) );
  NAND2_X1 U405 ( .A1(n351), .A2(n349), .ZN(G60) );
  NAND2_X1 U406 ( .A1(n359), .A2(n350), .ZN(n349) );
  AND2_X1 U407 ( .A1(n357), .A2(n363), .ZN(n350) );
  NOR2_X1 U408 ( .A1(n355), .A2(n352), .ZN(n351) );
  NAND2_X1 U409 ( .A1(n354), .A2(n353), .ZN(n352) );
  OR2_X1 U410 ( .A1(n357), .A2(n356), .ZN(n354) );
  NOR2_X1 U411 ( .A1(n359), .A2(n356), .ZN(n355) );
  NAND2_X1 U412 ( .A1(n742), .A2(n358), .ZN(n357) );
  NOR2_X1 U413 ( .A1(n365), .A2(n361), .ZN(n358) );
  NOR2_X1 U414 ( .A1(n362), .A2(n360), .ZN(n359) );
  INV_X1 U415 ( .A(G475), .ZN(n361) );
  INV_X1 U416 ( .A(KEYINPUT60), .ZN(n363) );
  INV_X1 U417 ( .A(n657), .ZN(n365) );
  XNOR2_X1 U418 ( .A(G902), .B(KEYINPUT15), .ZN(n638) );
  XNOR2_X1 U419 ( .A(n534), .B(KEYINPUT6), .ZN(n623) );
  XNOR2_X1 U420 ( .A(n766), .B(n472), .ZN(n485) );
  OR2_X1 U421 ( .A1(n534), .A2(n537), .ZN(n408) );
  XNOR2_X1 U422 ( .A(n613), .B(n422), .ZN(n615) );
  INV_X1 U423 ( .A(KEYINPUT47), .ZN(n422) );
  NAND2_X1 U424 ( .A1(n640), .A2(n637), .ZN(n456) );
  NOR2_X1 U425 ( .A1(n638), .A2(KEYINPUT65), .ZN(n455) );
  OR2_X1 U426 ( .A1(n366), .A2(n457), .ZN(n454) );
  INV_X1 U427 ( .A(G237), .ZN(n491) );
  INV_X1 U428 ( .A(KEYINPUT48), .ZN(n437) );
  XNOR2_X1 U429 ( .A(KEYINPUT70), .B(G137), .ZN(n470) );
  AND2_X1 U430 ( .A1(n380), .A2(n379), .ZN(n375) );
  NOR2_X1 U431 ( .A1(n382), .A2(n381), .ZN(n378) );
  AND2_X1 U432 ( .A1(n429), .A2(n428), .ZN(n427) );
  NAND2_X1 U433 ( .A1(G469), .A2(n426), .ZN(n425) );
  NOR2_X1 U434 ( .A1(n646), .A2(G902), .ZN(n396) );
  BUF_X1 U435 ( .A(n623), .Z(n400) );
  XNOR2_X1 U436 ( .A(n418), .B(n416), .ZN(n509) );
  XNOR2_X1 U437 ( .A(KEYINPUT86), .B(KEYINPUT8), .ZN(n418) );
  NOR2_X1 U438 ( .A1(n417), .A2(G953), .ZN(n416) );
  INV_X1 U439 ( .A(G234), .ZN(n417) );
  XNOR2_X1 U440 ( .A(n462), .B(n368), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n519), .B(KEYINPUT10), .ZN(n500) );
  NOR2_X2 U442 ( .A1(n701), .A2(n707), .ZN(n412) );
  XNOR2_X1 U443 ( .A(n593), .B(KEYINPUT39), .ZN(n436) );
  XNOR2_X1 U444 ( .A(n421), .B(n420), .ZN(n419) );
  INV_X1 U445 ( .A(KEYINPUT76), .ZN(n420) );
  XNOR2_X1 U446 ( .A(n690), .B(KEYINPUT89), .ZN(n438) );
  INV_X1 U447 ( .A(n597), .ZN(n382) );
  INV_X1 U448 ( .A(KEYINPUT78), .ZN(n381) );
  NAND2_X1 U449 ( .A1(n665), .A2(G902), .ZN(n428) );
  NOR2_X1 U450 ( .A1(G953), .A2(n732), .ZN(n481) );
  XNOR2_X1 U451 ( .A(n459), .B(KEYINPUT20), .ZN(n466) );
  NAND2_X1 U452 ( .A1(n366), .A2(KEYINPUT65), .ZN(n451) );
  NAND2_X1 U453 ( .A1(n454), .A2(n453), .ZN(n452) );
  NAND2_X1 U454 ( .A1(n366), .A2(n373), .ZN(n453) );
  XNOR2_X1 U455 ( .A(G116), .B(KEYINPUT5), .ZN(n488) );
  INV_X1 U456 ( .A(KEYINPUT68), .ZN(n404) );
  INV_X1 U457 ( .A(KEYINPUT75), .ZN(n431) );
  NOR2_X1 U458 ( .A1(G953), .A2(G237), .ZN(n495) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n524) );
  XNOR2_X1 U460 ( .A(n401), .B(n478), .ZN(n482) );
  XNOR2_X1 U461 ( .A(n402), .B(KEYINPUT14), .ZN(n401) );
  INV_X1 U462 ( .A(KEYINPUT77), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n444), .A2(n535), .ZN(n443) );
  NAND2_X1 U464 ( .A1(n466), .A2(G217), .ZN(n415) );
  XNOR2_X1 U465 ( .A(n391), .B(n437), .ZN(n636) );
  XOR2_X1 U466 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n506) );
  INV_X1 U467 ( .A(G134), .ZN(n469) );
  XNOR2_X1 U468 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n493) );
  XNOR2_X1 U469 ( .A(n485), .B(n477), .ZN(n667) );
  XNOR2_X1 U470 ( .A(n473), .B(KEYINPUT97), .ZN(n474) );
  NOR2_X1 U471 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U472 ( .A1(n619), .A2(n704), .ZN(n620) );
  BUF_X1 U473 ( .A(n714), .Z(n403) );
  INV_X1 U474 ( .A(KEYINPUT90), .ZN(n410) );
  INV_X2 U475 ( .A(G953), .ZN(n770) );
  XNOR2_X1 U476 ( .A(n461), .B(n465), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n384), .B(n500), .ZN(n383) );
  XNOR2_X1 U478 ( .A(n604), .B(KEYINPUT113), .ZN(n781) );
  AND2_X1 U479 ( .A1(n372), .A2(n456), .ZN(n366) );
  XOR2_X1 U480 ( .A(n490), .B(n407), .Z(n367) );
  INV_X1 U481 ( .A(KEYINPUT65), .ZN(n457) );
  XOR2_X1 U482 ( .A(G128), .B(G137), .Z(n368) );
  AND2_X1 U483 ( .A1(G214), .A2(n495), .ZN(n369) );
  AND2_X1 U484 ( .A1(n403), .A2(n596), .ZN(n371) );
  INV_X1 U485 ( .A(G902), .ZN(n426) );
  OR2_X1 U486 ( .A1(n640), .A2(n639), .ZN(n372) );
  OR2_X1 U487 ( .A1(n640), .A2(n457), .ZN(n373) );
  NAND2_X1 U488 ( .A1(n375), .A2(n377), .ZN(n374) );
  NAND2_X1 U489 ( .A1(n376), .A2(n378), .ZN(n377) );
  INV_X1 U490 ( .A(n572), .ZN(n376) );
  NAND2_X1 U491 ( .A1(n382), .A2(n381), .ZN(n379) );
  NAND2_X1 U492 ( .A1(n572), .A2(n381), .ZN(n380) );
  OR2_X1 U493 ( .A1(n667), .A2(n425), .ZN(n424) );
  INV_X1 U494 ( .A(n742), .ZN(n385) );
  BUF_X1 U495 ( .A(n659), .Z(n386) );
  INV_X1 U496 ( .A(n666), .ZN(n387) );
  AND2_X1 U497 ( .A1(n397), .A2(n580), .ZN(n399) );
  INV_X1 U498 ( .A(n666), .ZN(n742) );
  BUF_X1 U499 ( .A(n742), .Z(n747) );
  XNOR2_X2 U500 ( .A(n564), .B(n563), .ZN(n664) );
  AND2_X2 U501 ( .A1(n588), .A2(n654), .ZN(n565) );
  XNOR2_X1 U502 ( .A(n485), .B(n367), .ZN(n646) );
  BUF_X1 U503 ( .A(n397), .Z(n388) );
  XNOR2_X1 U504 ( .A(n586), .B(n585), .ZN(n397) );
  XNOR2_X2 U505 ( .A(n516), .B(n389), .ZN(n406) );
  XNOR2_X1 U506 ( .A(n389), .B(n489), .ZN(n407) );
  XNOR2_X2 U507 ( .A(n398), .B(G119), .ZN(n389) );
  NAND2_X1 U508 ( .A1(n705), .A2(n390), .ZN(n593) );
  NOR2_X2 U509 ( .A1(n778), .A2(n781), .ZN(n395) );
  NAND2_X1 U510 ( .A1(n390), .A2(n533), .ZN(n606) );
  NAND2_X1 U511 ( .A1(n394), .A2(n392), .ZN(n391) );
  XNOR2_X1 U512 ( .A(n393), .B(KEYINPUT71), .ZN(n392) );
  NAND2_X1 U513 ( .A1(n419), .A2(n438), .ZN(n393) );
  XNOR2_X1 U514 ( .A(n395), .B(KEYINPUT46), .ZN(n394) );
  XNOR2_X2 U515 ( .A(n396), .B(G472), .ZN(n534) );
  XNOR2_X1 U516 ( .A(n388), .B(n782), .ZN(G3) );
  XNOR2_X2 U517 ( .A(G113), .B(KEYINPUT3), .ZN(n398) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n430) );
  NAND2_X1 U519 ( .A1(n409), .A2(n371), .ZN(n586) );
  NAND2_X1 U520 ( .A1(n581), .A2(n399), .ZN(n435) );
  XNOR2_X1 U521 ( .A(n584), .B(n410), .ZN(n409) );
  AND2_X2 U522 ( .A1(n779), .A2(n664), .ZN(n589) );
  XNOR2_X1 U523 ( .A(n405), .B(n404), .ZN(n433) );
  XNOR2_X2 U524 ( .A(KEYINPUT67), .B(G101), .ZN(n471) );
  XNOR2_X2 U525 ( .A(n765), .B(n471), .ZN(n521) );
  XNOR2_X2 U526 ( .A(n406), .B(n518), .ZN(n759) );
  NAND2_X1 U527 ( .A1(n654), .A2(n587), .ZN(n405) );
  NAND2_X1 U528 ( .A1(n616), .A2(n617), .ZN(n421) );
  NAND2_X1 U529 ( .A1(n641), .A2(n455), .ZN(n450) );
  AND2_X2 U530 ( .A1(n752), .A2(n411), .ZN(n641) );
  INV_X1 U531 ( .A(n769), .ZN(n411) );
  XNOR2_X2 U532 ( .A(n414), .B(n345), .ZN(n596) );
  NOR2_X2 U533 ( .A1(n748), .A2(G902), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n667), .A2(n665), .ZN(n429) );
  NAND2_X2 U535 ( .A1(n427), .A2(n424), .ZN(n600) );
  NAND2_X1 U536 ( .A1(n434), .A2(n430), .ZN(n591) );
  NAND2_X1 U537 ( .A1(n433), .A2(n589), .ZN(n432) );
  XNOR2_X1 U538 ( .A(n435), .B(KEYINPUT91), .ZN(n434) );
  NAND2_X1 U539 ( .A1(n436), .A2(n592), .ZN(n595) );
  NAND2_X1 U540 ( .A1(n436), .A2(n687), .ZN(n692) );
  AND2_X2 U541 ( .A1(n583), .A2(n716), .ZN(n562) );
  NAND2_X2 U542 ( .A1(n642), .A2(n699), .ZN(n643) );
  XNOR2_X1 U543 ( .A(n439), .B(n519), .ZN(n520) );
  XNOR2_X2 U544 ( .A(n439), .B(n469), .ZN(n507) );
  XNOR2_X2 U545 ( .A(G143), .B(G128), .ZN(n439) );
  AND2_X1 U546 ( .A1(n441), .A2(n440), .ZN(n446) );
  NAND2_X1 U547 ( .A1(n714), .A2(n535), .ZN(n440) );
  NAND2_X1 U548 ( .A1(n442), .A2(n623), .ZN(n441) );
  NOR2_X1 U549 ( .A1(n714), .A2(n447), .ZN(n442) );
  NAND2_X1 U550 ( .A1(n623), .A2(n445), .ZN(n444) );
  INV_X1 U551 ( .A(n713), .ZN(n445) );
  OR2_X2 U552 ( .A1(n449), .A2(n448), .ZN(n642) );
  NOR2_X1 U553 ( .A1(n641), .A2(n451), .ZN(n448) );
  NAND2_X1 U554 ( .A1(n450), .A2(n452), .ZN(n449) );
  NAND2_X1 U555 ( .A1(n747), .A2(G478), .ZN(n745) );
  XNOR2_X2 U556 ( .A(n511), .B(n510), .ZN(n516) );
  XNOR2_X2 U557 ( .A(G122), .B(G116), .ZN(n511) );
  OR2_X1 U558 ( .A1(n713), .A2(n600), .ZN(n572) );
  XNOR2_X2 U559 ( .A(n630), .B(KEYINPUT38), .ZN(n705) );
  INV_X1 U560 ( .A(KEYINPUT84), .ZN(n607) );
  INV_X1 U561 ( .A(n618), .ZN(n619) );
  XNOR2_X1 U562 ( .A(n503), .B(G475), .ZN(n504) );
  INV_X1 U563 ( .A(n743), .ZN(n744) );
  XNOR2_X1 U564 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U565 ( .A1(G234), .A2(n638), .ZN(n459) );
  NAND2_X1 U566 ( .A1(G221), .A2(n466), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n460), .B(KEYINPUT21), .ZN(n717) );
  XNOR2_X1 U568 ( .A(n717), .B(KEYINPUT98), .ZN(n551) );
  INV_X1 U569 ( .A(n551), .ZN(n468) );
  XNOR2_X2 U570 ( .A(G146), .B(G125), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n509), .A2(G221), .ZN(n461) );
  XOR2_X1 U572 ( .A(G110), .B(G119), .Z(n462) );
  XOR2_X1 U573 ( .A(KEYINPUT73), .B(KEYINPUT23), .Z(n464) );
  XNOR2_X1 U574 ( .A(G140), .B(KEYINPUT24), .ZN(n463) );
  XNOR2_X1 U575 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U576 ( .A(KEYINPUT25), .B(KEYINPUT79), .ZN(n467) );
  NAND2_X1 U577 ( .A1(n468), .A2(n596), .ZN(n713) );
  XNOR2_X2 U578 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n765) );
  XNOR2_X1 U579 ( .A(n521), .B(G146), .ZN(n472) );
  XNOR2_X1 U580 ( .A(G107), .B(n501), .ZN(n475) );
  NAND2_X1 U581 ( .A1(n770), .A2(G227), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U583 ( .A(G110), .B(G104), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n476), .B(n517), .ZN(n477) );
  INV_X1 U585 ( .A(G469), .ZN(n665) );
  NAND2_X1 U586 ( .A1(G234), .A2(G237), .ZN(n478) );
  NAND2_X1 U587 ( .A1(n482), .A2(G952), .ZN(n479) );
  XOR2_X1 U588 ( .A(KEYINPUT95), .B(n479), .Z(n732) );
  INV_X1 U589 ( .A(KEYINPUT96), .ZN(n480) );
  XNOR2_X1 U590 ( .A(n481), .B(n480), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G902), .A2(n482), .ZN(n539) );
  NOR2_X1 U592 ( .A1(G900), .A2(n539), .ZN(n483) );
  NAND2_X1 U593 ( .A1(G953), .A2(n483), .ZN(n484) );
  NAND2_X1 U594 ( .A1(n542), .A2(n484), .ZN(n597) );
  XOR2_X1 U595 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n487) );
  NAND2_X1 U596 ( .A1(n495), .A2(G210), .ZN(n486) );
  XNOR2_X1 U597 ( .A(n487), .B(n486), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n488), .B(G131), .ZN(n489) );
  INV_X1 U599 ( .A(G472), .ZN(n644) );
  NAND2_X1 U600 ( .A1(n426), .A2(n491), .ZN(n528) );
  INV_X1 U601 ( .A(n704), .ZN(n537) );
  INV_X1 U602 ( .A(n492), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n496), .B(n369), .ZN(n499) );
  XNOR2_X1 U605 ( .A(n370), .B(n497), .ZN(n498) );
  XNOR2_X1 U606 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U607 ( .A(n501), .B(n500), .ZN(n767) );
  XNOR2_X1 U608 ( .A(n502), .B(n767), .ZN(n656) );
  INV_X1 U609 ( .A(KEYINPUT13), .ZN(n503) );
  XNOR2_X2 U610 ( .A(n505), .B(n504), .ZN(n576) );
  XNOR2_X1 U611 ( .A(n506), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U612 ( .A(n507), .B(n508), .ZN(n514) );
  NAND2_X1 U613 ( .A1(G217), .A2(n509), .ZN(n512) );
  INV_X1 U614 ( .A(G107), .ZN(n510) );
  XNOR2_X1 U615 ( .A(n516), .B(n512), .ZN(n513) );
  XNOR2_X1 U616 ( .A(n514), .B(n513), .ZN(n743) );
  NAND2_X1 U617 ( .A1(n743), .A2(n426), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n515), .B(G478), .ZN(n575) );
  INV_X1 U619 ( .A(n575), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n576), .A2(n550), .ZN(n546) );
  INV_X1 U621 ( .A(n546), .ZN(n532) );
  XNOR2_X1 U622 ( .A(n517), .B(KEYINPUT16), .ZN(n518) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n526) );
  NAND2_X1 U624 ( .A1(G224), .A2(n770), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n522), .B(KEYINPUT80), .ZN(n523) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n527), .B(n759), .ZN(n659) );
  INV_X1 U629 ( .A(n638), .ZN(n640) );
  NOR2_X1 U630 ( .A1(n659), .A2(n640), .ZN(n531) );
  NAND2_X1 U631 ( .A1(n528), .A2(G210), .ZN(n529) );
  XOR2_X1 U632 ( .A(n529), .B(KEYINPUT94), .Z(n530) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n536) );
  BUF_X2 U634 ( .A(n536), .Z(n630) );
  NOR2_X1 U635 ( .A1(n532), .A2(n630), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n606), .B(G143), .ZN(G45) );
  INV_X1 U637 ( .A(KEYINPUT63), .ZN(n653) );
  XNOR2_X1 U638 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n535) );
  INV_X1 U639 ( .A(n536), .ZN(n538) );
  INV_X1 U640 ( .A(n539), .ZN(n540) );
  NOR2_X1 U641 ( .A1(G898), .A2(n770), .ZN(n760) );
  NAND2_X1 U642 ( .A1(n540), .A2(n760), .ZN(n541) );
  NAND2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U644 ( .A(KEYINPUT0), .ZN(n544) );
  BUF_X2 U645 ( .A(n554), .Z(n574) );
  NAND2_X1 U646 ( .A1(n711), .A2(n574), .ZN(n545) );
  XNOR2_X1 U647 ( .A(n545), .B(n458), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U649 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n548) );
  XNOR2_X2 U650 ( .A(n549), .B(n548), .ZN(n654) );
  NOR2_X1 U651 ( .A1(n707), .A2(n551), .ZN(n552) );
  XNOR2_X1 U652 ( .A(n552), .B(KEYINPUT106), .ZN(n553) );
  NAND2_X1 U653 ( .A1(n554), .A2(n553), .ZN(n556) );
  INV_X1 U654 ( .A(KEYINPUT22), .ZN(n555) );
  XNOR2_X1 U655 ( .A(n556), .B(n555), .ZN(n583) );
  INV_X1 U656 ( .A(n596), .ZN(n716) );
  AND2_X1 U657 ( .A1(n403), .A2(n719), .ZN(n557) );
  NAND2_X1 U658 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X2 U659 ( .A(n558), .B(KEYINPUT108), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n400), .B(KEYINPUT83), .ZN(n560) );
  INV_X1 U661 ( .A(n403), .ZN(n559) );
  AND2_X1 U662 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U663 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U664 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n563) );
  NAND2_X1 U665 ( .A1(n565), .A2(n664), .ZN(n566) );
  NAND2_X1 U666 ( .A1(n566), .A2(KEYINPUT44), .ZN(n581) );
  OR2_X1 U667 ( .A1(n713), .A2(n719), .ZN(n567) );
  OR2_X1 U668 ( .A1(n403), .A2(n567), .ZN(n724) );
  INV_X1 U669 ( .A(n724), .ZN(n568) );
  NAND2_X1 U670 ( .A1(n574), .A2(n568), .ZN(n570) );
  XOR2_X1 U671 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n569) );
  XNOR2_X1 U672 ( .A(n570), .B(n569), .ZN(n688) );
  INV_X1 U673 ( .A(n719), .ZN(n571) );
  NOR2_X1 U674 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U675 ( .A1(n574), .A2(n573), .ZN(n677) );
  OR2_X1 U676 ( .A1(n688), .A2(n677), .ZN(n579) );
  AND2_X1 U677 ( .A1(n576), .A2(n575), .ZN(n687) );
  XNOR2_X2 U678 ( .A(KEYINPUT105), .B(n577), .ZN(n702) );
  INV_X1 U679 ( .A(n702), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U681 ( .A(n400), .ZN(n582) );
  NAND2_X1 U682 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U683 ( .A(KEYINPUT107), .ZN(n585) );
  INV_X1 U684 ( .A(KEYINPUT44), .ZN(n587) );
  BUF_X2 U685 ( .A(n588), .Z(n779) );
  XNOR2_X1 U686 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n590) );
  XNOR2_X1 U687 ( .A(n591), .B(n590), .ZN(n752) );
  XOR2_X1 U688 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n594) );
  XNOR2_X1 U689 ( .A(n595), .B(n594), .ZN(n778) );
  NOR2_X1 U690 ( .A1(n717), .A2(n596), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U692 ( .A(KEYINPUT72), .B(n599), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n600), .B(KEYINPUT111), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n612), .A2(n610), .ZN(n601) );
  NOR2_X1 U695 ( .A1(n601), .A2(n734), .ZN(n603) );
  INV_X1 U696 ( .A(KEYINPUT42), .ZN(n602) );
  XNOR2_X1 U697 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U698 ( .A1(n702), .A2(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U699 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U700 ( .A(n608), .B(n607), .ZN(n617) );
  AND2_X1 U701 ( .A1(n609), .A2(n610), .ZN(n611) );
  NAND2_X1 U702 ( .A1(n613), .A2(n702), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U704 ( .A(n592), .ZN(n621) );
  INV_X1 U705 ( .A(n630), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n627), .A2(n624), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n625), .B(KEYINPUT36), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n403), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n628) );
  XNOR2_X1 U710 ( .A(n629), .B(n628), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n633) );
  INV_X1 U712 ( .A(KEYINPUT110), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n633), .B(n632), .ZN(n780) );
  INV_X1 U714 ( .A(n780), .ZN(n634) );
  AND2_X1 U715 ( .A1(n634), .A2(n692), .ZN(n635) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n696) );
  NOR2_X1 U717 ( .A1(n696), .A2(KEYINPUT87), .ZN(n637) );
  NAND2_X1 U718 ( .A1(KEYINPUT2), .A2(KEYINPUT87), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n694), .A2(KEYINPUT2), .ZN(n699) );
  XNOR2_X2 U720 ( .A(n643), .B(KEYINPUT64), .ZN(n666) );
  NOR2_X1 U721 ( .A1(n666), .A2(n644), .ZN(n648) );
  XOR2_X1 U722 ( .A(KEYINPUT92), .B(KEYINPUT62), .Z(n645) );
  XNOR2_X1 U723 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n648), .B(n647), .ZN(n651) );
  INV_X1 U725 ( .A(G952), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n649), .A2(G953), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(G57) );
  BUF_X1 U728 ( .A(n654), .Z(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(G122), .ZN(G24) );
  XOR2_X1 U730 ( .A(KEYINPUT59), .B(n656), .Z(n657) );
  NAND2_X1 U731 ( .A1(n387), .A2(G210), .ZN(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  XNOR2_X1 U733 ( .A(n386), .B(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U735 ( .A1(n662), .A2(n751), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U737 ( .A(n664), .B(G119), .ZN(G21) );
  NOR2_X1 U738 ( .A1(n385), .A2(n665), .ZN(n671) );
  BUF_X1 U739 ( .A(n667), .Z(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n672), .A2(n751), .ZN(G54) );
  NAND2_X1 U744 ( .A1(n677), .A2(n592), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n673), .B(G104), .ZN(G6) );
  XOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n675) );
  XNOR2_X1 U747 ( .A(G107), .B(KEYINPUT115), .ZN(n674) );
  XNOR2_X1 U748 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U749 ( .A(KEYINPUT26), .B(n676), .Z(n679) );
  NAND2_X1 U750 ( .A1(n677), .A2(n687), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(G9) );
  XOR2_X1 U752 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U753 ( .A1(n613), .A2(n687), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U755 ( .A(G128), .B(n682), .Z(G30) );
  XOR2_X1 U756 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n684) );
  NAND2_X1 U757 ( .A1(n613), .A2(n592), .ZN(n683) );
  XNOR2_X1 U758 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U759 ( .A(G146), .B(n685), .ZN(G48) );
  NAND2_X1 U760 ( .A1(n592), .A2(n688), .ZN(n686) );
  XNOR2_X1 U761 ( .A(G113), .B(n686), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U763 ( .A(n689), .B(G116), .ZN(G18) );
  XNOR2_X1 U764 ( .A(G125), .B(n690), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n691), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U766 ( .A(G134), .B(KEYINPUT120), .ZN(n693) );
  XNOR2_X1 U767 ( .A(n693), .B(n692), .ZN(G36) );
  NOR2_X1 U768 ( .A1(n694), .A2(KEYINPUT85), .ZN(n695) );
  NOR2_X1 U769 ( .A1(n695), .A2(KEYINPUT2), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n696), .A2(KEYINPUT85), .ZN(n697) );
  OR2_X1 U771 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n738) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(n703), .Z(n710) );
  NOR2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(KEYINPUT122), .B(n708), .ZN(n709) );
  NOR2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n712) );
  INV_X1 U779 ( .A(n711), .ZN(n733) );
  NOR2_X1 U780 ( .A1(n712), .A2(n733), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n403), .A2(n713), .ZN(n715) );
  XNOR2_X1 U782 ( .A(n715), .B(KEYINPUT50), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U784 ( .A(KEYINPUT49), .B(n718), .Z(n720) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(n721), .B(KEYINPUT121), .ZN(n722) );
  NAND2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U789 ( .A(KEYINPUT51), .B(n726), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n727), .A2(n734), .ZN(n728) );
  NOR2_X1 U791 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT52), .ZN(n731) );
  NOR2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n736) );
  NOR2_X1 U794 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U795 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U796 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U797 ( .A(KEYINPUT124), .B(n739), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n740), .A2(G953), .ZN(n741) );
  XNOR2_X1 U799 ( .A(n741), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U800 ( .A1(n751), .A2(n746), .ZN(G63) );
  NAND2_X1 U801 ( .A1(n747), .A2(G217), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U803 ( .A1(n751), .A2(n750), .ZN(G66) );
  BUF_X1 U804 ( .A(n752), .Z(n753) );
  NAND2_X1 U805 ( .A1(n753), .A2(n770), .ZN(n754) );
  XOR2_X1 U806 ( .A(KEYINPUT125), .B(n754), .Z(n758) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n755), .ZN(n756) );
  NAND2_X1 U809 ( .A1(n756), .A2(G898), .ZN(n757) );
  NAND2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n763) );
  XOR2_X1 U811 ( .A(n759), .B(G101), .Z(n761) );
  NOR2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U814 ( .A(KEYINPUT126), .B(n764), .ZN(G69) );
  XNOR2_X1 U815 ( .A(n765), .B(n766), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(n772) );
  XNOR2_X1 U817 ( .A(n769), .B(n772), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(n770), .ZN(n777) );
  XNOR2_X1 U819 ( .A(G227), .B(n772), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U821 ( .A1(G953), .A2(n774), .ZN(n775) );
  XOR2_X1 U822 ( .A(KEYINPUT127), .B(n775), .Z(n776) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U824 ( .A(G131), .B(n778), .Z(G33) );
  XNOR2_X1 U825 ( .A(n779), .B(G110), .ZN(G12) );
  XOR2_X1 U826 ( .A(G140), .B(n780), .Z(G42) );
  XOR2_X1 U827 ( .A(n781), .B(G137), .Z(G39) );
  XNOR2_X1 U828 ( .A(G101), .B(KEYINPUT114), .ZN(n782) );
endmodule

