//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n215), .B1(new_n216), .B2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G13), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n218), .A2(KEYINPUT66), .A3(G1), .A4(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n214), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n213), .B1(new_n224), .B2(KEYINPUT0), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(KEYINPUT0), .B2(new_n224), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n223), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  INV_X1    g0033(.A(G97), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n232), .B1(new_n207), .B2(new_n233), .C1(new_n234), .C2(new_n222), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n216), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(new_n212), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n211), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n254), .A2(new_n212), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G50), .B1(new_n211), .B2(G1), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n269), .A2(new_n270), .B1(G50), .B2(new_n265), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G222), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(G1698), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT68), .B(G223), .Z(new_n281));
  OAI221_X1 g0081(.A(new_n279), .B1(new_n228), .B2(new_n277), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n289), .A3(G274), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT67), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(KEYINPUT67), .A3(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n291), .B1(new_n296), .B2(G226), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G179), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI211_X1 g0100(.A(new_n272), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n284), .A2(G190), .A3(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n298), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n260), .A2(G50), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT71), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n311), .B(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n259), .A2(G77), .B1(G20), .B2(new_n208), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n267), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT11), .B(new_n267), .C1(new_n313), .C2(new_n315), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT12), .B1(new_n265), .B2(G68), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n208), .B1(new_n264), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n321), .B1(new_n268), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT72), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  OAI211_X1 g0128(.A(G232), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(G226), .B(new_n278), .C1(new_n327), .C2(new_n328), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n283), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n289), .A2(KEYINPUT67), .A3(new_n292), .ZN(new_n334));
  OAI21_X1  g0134(.A(G238), .B1(new_n334), .B2(new_n293), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(new_n290), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT70), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n326), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT70), .A4(new_n290), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n333), .A2(new_n335), .A3(new_n326), .A4(new_n290), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G190), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G200), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n325), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT73), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n291), .B1(new_n296), .B2(G244), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n230), .C2(new_n277), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n283), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n300), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n257), .A2(new_n260), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n355), .B1(new_n211), .B2(new_n228), .C1(new_n258), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n267), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n228), .B1(new_n264), .B2(G20), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n268), .A2(new_n359), .B1(new_n228), .B2(new_n266), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n348), .A2(new_n362), .A3(new_n352), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n354), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n348), .B2(new_n352), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(KEYINPUT69), .B1(new_n353), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n348), .A2(G190), .A3(new_n352), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n346), .A2(KEYINPUT73), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n310), .A2(new_n347), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n256), .B1(new_n264), .B2(G20), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n268), .B1(new_n266), .B2(new_n256), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n327), .A2(new_n328), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n377), .B2(new_n211), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n276), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n202), .ZN(new_n384));
  INV_X1    g0184(.A(G159), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n385), .A2(G20), .A3(G33), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT75), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n211), .B1(new_n209), .B2(new_n382), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT75), .B1(new_n390), .B2(new_n386), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n267), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n275), .A2(new_n211), .A3(new_n276), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n379), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(G68), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n391), .A2(new_n389), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n376), .B1(new_n393), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(G223), .A2(G1698), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n404), .B1(G226), .B2(new_n278), .C1(new_n327), .C2(new_n328), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n283), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n289), .A2(new_n292), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n290), .B1(new_n233), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n300), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n289), .B1(new_n405), .B2(new_n406), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n413), .A2(new_n410), .A3(new_n362), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n403), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n408), .A2(new_n411), .A3(new_n367), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n365), .B1(new_n413), .B2(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n376), .B(new_n423), .C1(new_n393), .C2(new_n402), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n400), .A2(new_n401), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n391), .A2(new_n389), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n208), .B1(new_n396), .B2(new_n379), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n255), .B1(new_n432), .B2(KEYINPUT16), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n376), .A4(new_n423), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n418), .A2(new_n420), .A3(new_n426), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n341), .A2(G179), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n338), .B2(new_n339), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n344), .A2(G169), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n344), .A2(KEYINPUT74), .A3(KEYINPUT14), .A4(G169), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n325), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n374), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT78), .B1(new_n274), .B2(G1), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n264), .A3(G33), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n268), .A2(G116), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT81), .B(G116), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n266), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n267), .B1(new_n460), .B2(new_n211), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n211), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n234), .A2(KEYINPUT77), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G97), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n274), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n455), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n255), .B1(G20), .B2(new_n452), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT77), .B(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n211), .B(new_n462), .C1(new_n471), .C2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n454), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G264), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n278), .C1(new_n327), .C2(new_n328), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n277), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n283), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n264), .B(G45), .C1(new_n285), .C2(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT79), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n264), .A4(G45), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G270), .A3(new_n289), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n480), .A2(KEYINPUT79), .B1(KEYINPUT5), .B2(new_n285), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(G274), .A3(new_n289), .A4(new_n485), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n479), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n474), .A2(new_n491), .A3(new_n362), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(G200), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n474), .C1(new_n367), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n469), .A2(new_n473), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n451), .A2(new_n453), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n300), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n498), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n498), .B2(new_n491), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n493), .B(new_n495), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n283), .B1(new_n489), .B2(new_n485), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n504));
  OAI211_X1 g0304(.A(G250), .B(new_n278), .C1(new_n327), .C2(new_n328), .ZN(new_n505));
  INV_X1    g0305(.A(G294), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n274), .C2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(G264), .B1(new_n507), .B2(new_n283), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n367), .A3(new_n490), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n487), .A2(G264), .A3(new_n289), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n490), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n365), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n211), .B1(new_n327), .B2(new_n328), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(KEYINPUT84), .B2(KEYINPUT22), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n277), .A2(new_n520), .A3(new_n211), .A4(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n211), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n460), .A2(new_n211), .A3(G33), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n519), .A2(new_n522), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT24), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n527), .A2(new_n526), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n522), .A4(new_n519), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n267), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n268), .A2(new_n450), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n265), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n514), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n508), .A2(new_n362), .A3(new_n490), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n512), .A2(new_n300), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n255), .B1(new_n529), .B2(new_n532), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n502), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  AND2_X1   g0349(.A1(KEYINPUT4), .A2(G244), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n278), .B(new_n550), .C1(new_n327), .C2(new_n328), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n229), .B1(new_n275), .B2(new_n276), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n462), .C1(new_n552), .C2(KEYINPUT4), .ZN(new_n553));
  OAI21_X1  g0353(.A(G250), .B1(new_n327), .B2(new_n328), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n278), .B1(new_n554), .B2(KEYINPUT4), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n283), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n487), .A2(G257), .A3(new_n289), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n490), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n300), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n556), .A2(new_n362), .A3(new_n490), .A4(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n265), .A2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n535), .B2(new_n234), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n398), .A2(G107), .A3(new_n399), .ZN(new_n565));
  XOR2_X1   g0365(.A(G97), .B(G107), .Z(new_n566));
  NAND2_X1  g0366(.A1(new_n230), .A2(KEYINPUT6), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n566), .A2(KEYINPUT6), .B1(new_n471), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n564), .B1(new_n570), .B2(new_n267), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n549), .B1(new_n561), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n267), .ZN(new_n573));
  INV_X1    g0373(.A(new_n564), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(KEYINPUT80), .A3(new_n560), .A4(new_n559), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n558), .A2(G200), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n577), .C1(new_n367), .C2(new_n558), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n580));
  OAI211_X1 g0380(.A(G238), .B(new_n278), .C1(new_n327), .C2(new_n328), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n274), .C2(new_n452), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n283), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n214), .B1(new_n286), .B2(G1), .ZN(new_n584));
  INV_X1    g0384(.A(G274), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n264), .A2(new_n585), .A3(G45), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n289), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n300), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n587), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n362), .B(new_n589), .C1(new_n582), .C2(new_n283), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT82), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(G179), .A3(new_n587), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n589), .B1(new_n582), .B2(new_n283), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n593), .C1(new_n300), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n211), .B1(new_n331), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n518), .A2(new_n230), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n467), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n471), .B2(new_n258), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n277), .A2(new_n211), .A3(G68), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n267), .B1(new_n266), .B2(new_n356), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n535), .B2(new_n356), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n591), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n583), .A2(G190), .A3(new_n587), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n536), .A2(G87), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n606), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n594), .A2(new_n365), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n548), .A2(new_n579), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n446), .A2(new_n613), .ZN(G372));
  AND2_X1   g0414(.A1(new_n418), .A2(new_n420), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n444), .B1(new_n364), .B2(new_n346), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n435), .A2(new_n426), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n308), .A2(new_n309), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n301), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n592), .B1(new_n300), .B2(new_n594), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n604), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n546), .B(new_n493), .C1(new_n500), .C2(new_n501), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n608), .A2(new_n609), .B1(new_n621), .B2(new_n604), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n542), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n561), .A2(new_n571), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT26), .B1(new_n628), .B2(new_n624), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n611), .B1(new_n572), .B2(new_n576), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n620), .B1(new_n446), .B2(new_n633), .ZN(G369));
  NAND2_X1  g0434(.A1(new_n496), .A2(new_n497), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G169), .A3(new_n491), .ZN(new_n636));
  INV_X1    g0436(.A(new_n499), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n498), .A2(new_n491), .A3(new_n499), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n492), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n264), .A2(new_n211), .A3(G13), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n641), .A2(KEYINPUT85), .A3(KEYINPUT27), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT85), .B1(new_n641), .B2(KEYINPUT27), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(G213), .B1(new_n641), .B2(KEYINPUT27), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G343), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n547), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n546), .B2(new_n648), .ZN(new_n652));
  XOR2_X1   g0452(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  INV_X1    g0453(.A(new_n640), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n474), .A2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n502), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n534), .A2(new_n541), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n650), .B1(new_n661), .B2(new_n647), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n546), .B2(new_n647), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT87), .Z(G399));
  NOR3_X1   g0466(.A1(new_n221), .A2(KEYINPUT88), .A3(G41), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n220), .B2(new_n285), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n467), .A2(G116), .A3(new_n598), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n210), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n670), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT28), .Z(new_n676));
  INV_X1    g0476(.A(KEYINPUT29), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n677), .B(new_n647), .C1(new_n627), .C2(new_n631), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n624), .A2(new_n542), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n546), .B2(new_n640), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n680), .A2(new_n579), .B1(new_n621), .B2(new_n604), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n628), .B2(new_n624), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n630), .B2(new_n682), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n648), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n678), .B1(new_n685), .B2(new_n677), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n548), .A2(new_n579), .A3(new_n612), .A4(new_n647), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n590), .A2(new_n556), .A3(new_n490), .A4(new_n557), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n508), .A2(new_n490), .A3(new_n488), .A4(new_n479), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n558), .A2(new_n592), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n510), .A2(new_n511), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n491), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n594), .A2(G179), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n558), .A2(new_n697), .A3(new_n512), .A4(new_n491), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT31), .B1(new_n699), .B2(new_n648), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n687), .B1(new_n688), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n686), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n676), .B1(new_n704), .B2(G1), .ZN(G364));
  NOR2_X1   g0505(.A1(new_n218), .A2(G20), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n264), .B1(new_n706), .B2(G45), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n671), .A2(new_n707), .ZN(new_n708));
  OR3_X1    g0508(.A1(KEYINPUT91), .A2(G13), .A3(G33), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT91), .B1(G13), .B2(G33), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n212), .B1(G20), .B2(new_n300), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n249), .A2(new_n286), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n220), .A2(new_n377), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT89), .Z(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n286), .B2(new_n674), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n717), .B1(new_n722), .B2(KEYINPUT90), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(KEYINPUT90), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n221), .A2(new_n377), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(G355), .B1(new_n456), .B2(new_n221), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n716), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n211), .A2(new_n362), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(new_n367), .A3(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n211), .A2(G190), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n362), .A3(new_n365), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n730), .A2(G322), .B1(G329), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G311), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n734), .B(new_n377), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n362), .A2(G200), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n211), .A3(G190), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n738), .B1(G283), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n728), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(G317), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n367), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n211), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n743), .A2(new_n367), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G294), .A2(new_n751), .B1(new_n752), .B2(G326), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n742), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n740), .A2(new_n211), .A3(new_n367), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n754), .B1(G303), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n741), .A2(G107), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n756), .B2(new_n518), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n750), .A2(new_n234), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(G50), .B2(new_n752), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n377), .B1(new_n730), .B2(G58), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n765), .B(new_n766), .C1(new_n228), .C2(new_n737), .ZN(new_n767));
  OR3_X1    g0567(.A1(new_n732), .A2(KEYINPUT32), .A3(new_n385), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT32), .B1(new_n732), .B2(new_n385), .ZN(new_n769));
  INV_X1    g0569(.A(new_n744), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n208), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n763), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n761), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n708), .B(new_n727), .C1(new_n714), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n713), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n657), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n708), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n659), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G330), .B2(new_n657), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n364), .A2(new_n647), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n647), .B1(new_n358), .B2(new_n360), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n371), .B2(new_n368), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n784), .B2(new_n364), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n633), .B2(new_n648), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n372), .B(new_n647), .C1(new_n627), .C2(new_n631), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n688), .A2(new_n702), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G330), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n777), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n790), .B2(new_n788), .ZN(new_n792));
  INV_X1    g0592(.A(new_n714), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n712), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n777), .B1(G77), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n785), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n759), .A2(new_n230), .ZN(new_n798));
  INV_X1    g0598(.A(new_n741), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n518), .ZN(new_n800));
  INV_X1    g0600(.A(new_n730), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n377), .B1(new_n732), .B2(new_n735), .C1(new_n801), .C2(new_n506), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n798), .A2(new_n764), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n460), .A2(new_n736), .B1(new_n744), .B2(G283), .ZN(new_n804));
  INV_X1    g0604(.A(new_n752), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n477), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT94), .Z(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n730), .B1(new_n736), .B2(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G150), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n805), .C1(new_n810), .C2(new_n770), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n741), .A2(G68), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n377), .B1(new_n733), .B2(G132), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n207), .C2(new_n750), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n760), .B2(G50), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n803), .A2(new_n807), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n796), .B1(new_n797), .B2(new_n712), .C1(new_n793), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n792), .A2(new_n819), .ZN(G384));
  NOR2_X1   g0620(.A1(new_n706), .A2(new_n264), .ZN(new_n821));
  INV_X1    g0621(.A(new_n376), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n429), .B2(new_n433), .ZN(new_n823));
  INV_X1    g0623(.A(new_n646), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n435), .A2(new_n426), .A3(KEYINPUT100), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n418), .A3(new_n420), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT100), .B1(new_n435), .B2(new_n426), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n424), .B1(new_n823), .B2(new_n415), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT37), .B1(new_n830), .B2(new_n825), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n403), .A2(new_n646), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n417), .A2(new_n832), .A3(new_n833), .A4(new_n424), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n831), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n829), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n392), .A3(new_n267), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n824), .B1(new_n843), .B2(new_n376), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n436), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n424), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n415), .A2(new_n824), .B1(new_n843), .B2(new_n376), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n834), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n325), .A2(new_n342), .A3(new_n345), .ZN(new_n852));
  INV_X1    g0652(.A(new_n438), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n647), .A2(KEYINPUT73), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n344), .A2(G169), .B1(KEYINPUT74), .B2(KEYINPUT14), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n300), .B(new_n440), .C1(new_n343), .C2(new_n341), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n443), .B2(new_n648), .ZN(new_n858));
  INV_X1    g0658(.A(new_n325), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n852), .B(new_n785), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n789), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n851), .A2(KEYINPUT101), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n839), .B2(new_n840), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n789), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n845), .B2(new_n849), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n789), .A2(new_n797), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n445), .A2(new_n789), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n687), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n872), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n787), .B2(new_n782), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n870), .B2(new_n864), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n615), .A2(new_n646), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(KEYINPUT98), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n845), .A2(new_n849), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n840), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n850), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n850), .A2(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n841), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n443), .A2(new_n325), .A3(new_n648), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n885), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT98), .B1(new_n883), .B2(new_n884), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n686), .A2(new_n445), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n620), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  AOI21_X1  g0700(.A(new_n821), .B1(new_n880), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n880), .B2(new_n900), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n674), .A2(G77), .A3(new_n382), .ZN(new_n903));
  INV_X1    g0703(.A(new_n201), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n208), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G1), .A3(new_n218), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n212), .A2(new_n211), .A3(new_n456), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n568), .B2(KEYINPUT35), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT96), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n902), .A2(new_n906), .A3(new_n914), .ZN(G367));
  INV_X1    g0715(.A(new_n664), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n579), .B1(new_n571), .B2(new_n647), .ZN(new_n917));
  INV_X1    g0717(.A(new_n628), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n647), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT104), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n647), .B1(new_n603), .B2(new_n607), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT103), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n622), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n624), .B2(new_n923), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n921), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n919), .A2(new_n650), .A3(new_n649), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT42), .Z(new_n931));
  INV_X1    g0731(.A(new_n546), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n572), .A2(new_n576), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n647), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n929), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n928), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n670), .B(KEYINPUT41), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n653), .A2(new_n919), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n653), .A2(new_n919), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n653), .A2(new_n943), .A3(new_n919), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT45), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n946), .A2(new_n916), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n663), .A2(new_n649), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT106), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(KEYINPUT106), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n651), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n658), .ZN(new_n953));
  INV_X1    g0753(.A(new_n704), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n916), .B1(new_n946), .B2(new_n947), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n938), .B1(new_n957), .B2(new_n704), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n707), .B(KEYINPUT107), .Z(new_n959));
  OAI21_X1  g0759(.A(new_n937), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n720), .A2(new_n245), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n715), .B1(new_n220), .B2(new_n356), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n777), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n799), .A2(new_n228), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n377), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n751), .A2(G68), .ZN(new_n967));
  INV_X1    g0767(.A(G143), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(new_n770), .B2(new_n385), .C1(new_n968), .C2(new_n805), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n736), .A2(new_n904), .B1(G137), .B2(new_n733), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n810), .B2(new_n801), .C1(new_n756), .C2(new_n207), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n966), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(KEYINPUT108), .B2(new_n965), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT46), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n759), .A2(new_n974), .A3(new_n456), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n277), .B1(new_n733), .B2(G317), .ZN(new_n976));
  INV_X1    g0776(.A(G283), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(new_n737), .B2(new_n977), .C1(new_n477), .C2(new_n801), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n467), .B2(new_n741), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n974), .B1(new_n756), .B2(new_n452), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n770), .A2(new_n506), .B1(new_n805), .B2(new_n735), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G107), .B2(new_n751), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n973), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n963), .B1(new_n985), .B2(new_n714), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n925), .A2(new_n713), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n960), .A2(new_n988), .ZN(G387));
  INV_X1    g0789(.A(new_n955), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n953), .A2(new_n954), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n670), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n959), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n663), .A2(new_n775), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n719), .B1(new_n242), .B2(new_n286), .ZN(new_n995));
  INV_X1    g0795(.A(new_n725), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n672), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(G45), .B1(G68), .B2(G77), .ZN(new_n998));
  INV_X1    g0798(.A(G50), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n257), .A2(KEYINPUT50), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT50), .B1(new_n257), .B2(new_n999), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n672), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n997), .A2(new_n1002), .B1(new_n230), .B2(new_n221), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G303), .A2(new_n736), .B1(new_n730), .B2(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n735), .B2(new_n770), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G322), .B2(new_n752), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n756), .A2(new_n506), .B1(new_n977), .B2(new_n750), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT109), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(KEYINPUT109), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n799), .A2(new_n452), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n277), .B(new_n1014), .C1(G326), .C2(new_n733), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n377), .B1(new_n733), .B2(G150), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n737), .B2(new_n208), .C1(new_n999), .C2(new_n801), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n741), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n750), .A2(new_n356), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n770), .A2(new_n256), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G159), .C2(new_n752), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n755), .A2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n777), .B1(new_n716), .B2(new_n1003), .C1(new_n1025), .C2(new_n793), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n992), .B1(new_n953), .B2(new_n993), .C1(new_n994), .C2(new_n1026), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n948), .A2(new_n956), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT110), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n993), .B1(new_n1028), .B2(KEYINPUT110), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n919), .A2(new_n775), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n720), .A2(new_n252), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n715), .B1(new_n220), .B2(new_n471), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n777), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n750), .A2(new_n228), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n277), .B1(new_n968), .B2(new_n732), .C1(new_n737), .C2(new_n256), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n904), .C2(new_n744), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n208), .B2(new_n756), .C1(new_n518), .C2(new_n799), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n730), .A2(G159), .B1(new_n752), .B2(G150), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n730), .A2(G311), .B1(new_n752), .B2(G317), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n770), .A2(new_n477), .B1(new_n452), .B2(new_n750), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n377), .B1(new_n737), .B2(new_n506), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G322), .C2(new_n733), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n762), .C1(new_n977), .C2(new_n756), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1038), .A2(new_n1040), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1034), .B1(new_n1049), .B2(new_n714), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1028), .A2(new_n990), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n670), .A3(new_n957), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(G390));
  NAND2_X1  g0854(.A1(new_n841), .A2(new_n891), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT39), .B1(new_n864), .B2(new_n870), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n882), .C2(new_n893), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n703), .A2(new_n860), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n784), .A2(new_n364), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n934), .A2(new_n612), .A3(new_n682), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n683), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n647), .B(new_n1059), .C1(new_n627), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n782), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n872), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n851), .A3(new_n894), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1057), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n703), .A2(new_n860), .A3(KEYINPUT113), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n959), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n777), .B1(new_n257), .B2(new_n794), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n730), .A2(G132), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT54), .B(G143), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n277), .B1(new_n737), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G125), .C2(new_n733), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n770), .A2(new_n809), .B1(new_n385), .B2(new_n750), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G128), .B2(new_n752), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n201), .C2(new_n799), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n755), .A2(G150), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n759), .A2(new_n518), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n770), .A2(new_n230), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1035), .B(new_n1086), .C1(G283), .C2(new_n752), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n277), .B1(new_n733), .B2(G294), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n467), .A2(new_n736), .B1(new_n730), .B2(G116), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1087), .A2(new_n814), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1082), .A2(new_n1084), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1075), .B1(new_n1091), .B2(new_n714), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n838), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n837), .B1(new_n831), .B2(new_n834), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT38), .B1(new_n1095), .B2(new_n829), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1056), .B1(new_n1096), .B2(new_n890), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1097), .B2(new_n712), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n445), .A2(new_n703), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n898), .A2(new_n620), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n881), .B1(new_n790), .B2(new_n785), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n703), .A2(new_n860), .A3(KEYINPUT113), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT113), .B1(new_n703), .B2(new_n860), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n787), .A2(new_n782), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n789), .A2(KEYINPUT114), .A3(G330), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n797), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n703), .A2(KEYINPUT114), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n881), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1058), .A2(new_n782), .A3(new_n1063), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1102), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1100), .B1(new_n1073), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1057), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n787), .A2(new_n782), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n894), .B1(new_n1119), .B2(new_n881), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n865), .A2(new_n893), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1120), .A2(new_n892), .B1(new_n1121), .B2(new_n1065), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1118), .B1(new_n1122), .B2(new_n1071), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1102), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1071), .B2(new_n1103), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n785), .B1(new_n703), .B2(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(KEYINPUT114), .B2(new_n703), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1113), .B1(new_n1127), .B2(new_n881), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1124), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(KEYINPUT116), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1117), .A2(new_n670), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT115), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1071), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n893), .B1(new_n1107), .B2(new_n872), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1097), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n881), .B1(new_n1063), .B2(new_n782), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1136), .A2(new_n865), .A3(new_n893), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT115), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1116), .A2(new_n1138), .A3(new_n1139), .A4(new_n1118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1132), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1099), .B1(new_n1131), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1130), .A2(new_n670), .ZN(new_n1143));
  AND4_X1   g0943(.A1(new_n1099), .A2(new_n1143), .A3(new_n1141), .A4(new_n1117), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1074), .B(new_n1098), .C1(new_n1142), .C2(new_n1144), .ZN(G378));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1073), .B2(new_n1116), .ZN(new_n1146));
  AND4_X1   g0946(.A1(new_n1139), .A2(new_n1116), .A3(new_n1138), .A4(new_n1118), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1124), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n874), .A2(G330), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n868), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT120), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1149), .B1(new_n867), .B2(new_n862), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n272), .A2(new_n824), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT55), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n310), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1159));
  XOR2_X1   g0959(.A(new_n1158), .B(new_n1159), .Z(new_n1160));
  NAND3_X1  g0960(.A1(new_n1153), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1154), .A2(KEYINPUT120), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n897), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n897), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1154), .B2(KEYINPUT120), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n868), .A2(KEYINPUT120), .A3(new_n1150), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1163), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1165), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1148), .A2(KEYINPUT57), .A3(new_n1164), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT121), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1164), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1102), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1161), .A2(new_n897), .A3(new_n1163), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n897), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1141), .B2(new_n1124), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1172), .A2(new_n670), .A3(new_n1176), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1162), .A2(new_n711), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n777), .B1(new_n904), .B2(new_n794), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n967), .B1(new_n770), .B2(new_n234), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n741), .A2(G58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n377), .A2(new_n285), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n730), .B2(G107), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n356), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n736), .A2(new_n1190), .B1(G283), .B2(new_n733), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1023), .A2(new_n1187), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1186), .B(new_n1192), .C1(G116), .C2(new_n752), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1188), .B(new_n999), .C1(G33), .C2(G41), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n730), .A2(G128), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n737), .B2(new_n809), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G150), .B2(new_n751), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G125), .A2(new_n752), .B1(new_n744), .B2(G132), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n756), .C2(new_n1077), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n741), .A2(G159), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1197), .B1(KEYINPUT58), .B2(new_n1193), .C1(new_n1203), .C2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1208), .B2(new_n714), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1179), .A2(new_n959), .B1(new_n1184), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1183), .A2(new_n1210), .ZN(G375));
  OAI21_X1  g1011(.A(new_n959), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n881), .A2(new_n711), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n777), .B1(G68), .B2(new_n794), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n770), .A2(new_n1077), .B1(new_n999), .B2(new_n750), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G132), .B2(new_n752), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n377), .B1(new_n730), .B2(G137), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n736), .A2(G150), .B1(G128), .B2(new_n733), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1187), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(new_n759), .C2(new_n385), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1020), .B1(G283), .B2(new_n730), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT123), .Z(new_n1223));
  OAI221_X1 g1023(.A(new_n377), .B1(new_n477), .B2(new_n732), .C1(new_n737), .C2(new_n230), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n506), .A2(new_n805), .B1(new_n770), .B2(new_n452), .ZN(new_n1225));
  OR4_X1    g1025(.A1(new_n964), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n759), .A2(new_n234), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n1228), .B2(new_n714), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1212), .A2(KEYINPUT122), .B1(new_n1214), .B2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1213), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n938), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1108), .A2(new_n1115), .A3(new_n1102), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1129), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(G381));
  NOR2_X1   g1035(.A1(G390), .A2(G387), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1183), .A2(new_n1210), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1074), .A2(new_n1098), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1131), .B2(new_n1141), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .A4(new_n1240), .ZN(G407));
  INV_X1    g1041(.A(G213), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G343), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(new_n1239), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  NAND3_X1  g1045(.A1(new_n1183), .A2(G378), .A3(new_n1210), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1210), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1174), .A2(new_n938), .A3(new_n1175), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1239), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1243), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1233), .B(KEYINPUT60), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n670), .A3(new_n1129), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1231), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n792), .A3(new_n819), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1231), .A3(G384), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1253), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1243), .A2(G2897), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1260), .A2(new_n1253), .A3(new_n1262), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1250), .A2(new_n1251), .A3(new_n1260), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1243), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1272), .B2(new_n1260), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1267), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT127), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n780), .ZN(new_n1276));
  AND2_X1   g1076(.A1(G390), .A2(G387), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(new_n1236), .ZN(new_n1278));
  OR2_X1    g1078(.A1(G390), .A2(G387), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G390), .A2(G387), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1267), .B(new_n1284), .C1(new_n1271), .C2(new_n1273), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1275), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1272), .A2(new_n1260), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1283), .B1(KEYINPUT63), .B2(new_n1288), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(KEYINPUT124), .A3(KEYINPUT63), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1287), .B2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1267), .C1(new_n1290), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1286), .A2(new_n1294), .ZN(G405));
  AND2_X1   g1095(.A1(G375), .A2(new_n1239), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1246), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1260), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1298), .B(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1283), .ZN(G402));
endmodule


