//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  OR2_X1    g000(.A1(KEYINPUT65), .A2(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT65), .A2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G143), .ZN(new_n190));
  AOI22_X1  g004(.A1(G143), .A2(new_n189), .B1(new_n190), .B2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT0), .A3(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT64), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n187), .A2(new_n197), .A3(new_n188), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n192), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(new_n188), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(G143), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT64), .B(G143), .Z(new_n210));
  OAI211_X1 g024(.A(new_n207), .B(new_n209), .C1(new_n210), .C2(new_n194), .ZN(new_n211));
  INV_X1    g025(.A(new_n199), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT84), .B(G224), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n218), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n204), .A2(new_n221), .A3(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT6), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT76), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n234), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT77), .B(G101), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n230), .A2(G104), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n227), .A2(G107), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n233), .B2(new_n238), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT78), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n248), .B(new_n251), .C1(new_n233), .C2(new_n238), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n242), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n243), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n257), .A2(KEYINPUT5), .A3(G119), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(G113), .B2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n241), .A2(new_n245), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(G110), .B(G122), .Z(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n226), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n261), .A2(new_n263), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n261), .A2(new_n263), .A3(new_n226), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n224), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT7), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n221), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n220), .A2(new_n222), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n263), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n254), .A2(new_n260), .ZN(new_n274));
  INV_X1    g088(.A(new_n249), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n260), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n262), .B(KEYINPUT8), .Z(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n204), .A2(new_n270), .A3(new_n221), .A4(new_n216), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n272), .A2(new_n273), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(new_n269), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n268), .A2(new_n269), .A3(new_n282), .A4(new_n280), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT85), .A3(new_n285), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n281), .A2(KEYINPUT85), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT9), .B(G234), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n197), .B1(new_n187), .B2(new_n188), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  OAI21_X1  g113(.A(G128), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n199), .A2(new_n300), .B1(new_n191), .B2(new_n209), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n208), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n211), .B1(new_n191), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n253), .A2(new_n301), .B1(new_n275), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n305));
  INV_X1    g119(.A(G134), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G137), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(KEYINPUT11), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(G137), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT11), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT66), .B(new_n311), .C1(new_n306), .C2(G137), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n297), .B1(new_n304), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n253), .A2(new_n301), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n303), .A2(new_n275), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n316), .A2(KEYINPUT80), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(KEYINPUT80), .A3(new_n321), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n296), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n241), .A2(new_n203), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n254), .A2(KEYINPUT10), .A3(new_n214), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n308), .A2(new_n309), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n314), .A3(new_n310), .A4(new_n312), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n313), .A2(G131), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G140), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n218), .A2(G227), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n214), .B1(new_n250), .B2(new_n252), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n303), .A2(new_n275), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n334), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(new_n297), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n320), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT81), .B(new_n323), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n325), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT82), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n330), .A2(new_n334), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n339), .B1(new_n350), .B2(new_n335), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n325), .A2(new_n347), .A3(new_n352), .A4(new_n340), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G469), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n269), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n350), .A2(new_n335), .A3(new_n339), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n330), .A2(new_n334), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n322), .B2(new_n324), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n359), .B2(new_n339), .ZN(new_n360));
  OAI21_X1  g174(.A(G469), .B1(new_n360), .B2(G902), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n295), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n218), .A3(G214), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n210), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n364), .A2(G143), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT86), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT18), .A2(G131), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n367), .B(new_n368), .Z(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n189), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT73), .A2(G125), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(G140), .Z(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n373), .B2(new_n194), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n370), .A2(KEYINPUT19), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n373), .B2(KEYINPUT19), .ZN(new_n377));
  INV_X1    g191(.A(new_n189), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT88), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n365), .A2(new_n366), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n314), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n215), .A2(KEYINPUT16), .A3(G140), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G146), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n314), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n365), .A2(G131), .A3(new_n366), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(new_n383), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n379), .A2(KEYINPUT88), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n375), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(G113), .B(G122), .Z(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT89), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n227), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n385), .B(G146), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .A4(new_n366), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n389), .A2(new_n383), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(KEYINPUT17), .ZN(new_n401));
  INV_X1    g215(.A(new_n395), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n375), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n269), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT20), .ZN(new_n407));
  AOI21_X1  g221(.A(G475), .B1(new_n396), .B2(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n269), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n403), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n402), .B1(new_n401), .B2(new_n375), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n269), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G475), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G217), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n293), .A2(new_n417), .A3(G953), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n257), .A2(G122), .ZN(new_n419));
  INV_X1    g233(.A(G122), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n230), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT91), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n208), .A2(G143), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n210), .B2(new_n208), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(G134), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n421), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(KEYINPUT14), .B2(new_n419), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n424), .B(new_n427), .C1(new_n230), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n422), .B(G107), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n426), .A2(G134), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT13), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n190), .A2(new_n436), .A3(G128), .ZN(new_n437));
  OAI211_X1 g251(.A(G134), .B(new_n437), .C1(new_n426), .C2(new_n436), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n435), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n418), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n431), .A2(new_n440), .A3(new_n418), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G478), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(KEYINPUT93), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n443), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT93), .B(new_n269), .C1(new_n453), .C2(new_n441), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G952), .ZN(new_n457));
  AOI211_X1 g271(.A(G953), .B(new_n457), .C1(G234), .C2(G237), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(G898), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT94), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n269), .B(new_n218), .C1(G234), .C2(G237), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n416), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n291), .A2(new_n362), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G472), .ZN(new_n466));
  INV_X1    g280(.A(new_n310), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n467), .B2(new_n307), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n214), .A2(new_n332), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n192), .A2(new_n202), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n469), .B(new_n244), .C1(new_n315), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n203), .A2(new_n334), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n244), .B1(new_n474), .B2(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n474), .A2(new_n477), .A3(new_n244), .A4(new_n469), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n479), .B2(new_n472), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n363), .A2(new_n218), .A3(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G101), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n478), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n315), .A2(new_n470), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n214), .A2(new_n332), .A3(new_n468), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n474), .A2(KEYINPUT30), .A3(new_n469), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n245), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT29), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g311(.A(new_n485), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n479), .B2(new_n472), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(KEYINPUT29), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n466), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n487), .A2(new_n493), .A3(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n487), .A2(new_n493), .A3(KEYINPUT31), .A4(new_n498), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n480), .A2(new_n485), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G472), .A2(G902), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT69), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(KEYINPUT32), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n505), .A2(new_n506), .B1(new_n480), .B2(new_n485), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n511), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n509), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n512), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n502), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n417), .B1(G234), .B2(new_n269), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  XNOR2_X1  g336(.A(G119), .B(G128), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G110), .ZN(new_n525));
  OR2_X1    g339(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(G119), .A3(new_n208), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n523), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n397), .B(new_n524), .C1(new_n525), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n530), .A2(new_n532), .A3(new_n525), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n530), .B2(new_n525), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n522), .A2(new_n523), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n386), .A2(new_n371), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n531), .B(new_n541), .C1(new_n536), .C2(new_n537), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n269), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n521), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n544), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n521), .A2(G902), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n520), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n465), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n238), .ZN(G3));
  NOR2_X1   g372(.A1(new_n515), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n560));
  OAI21_X1  g374(.A(G472), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n509), .A2(new_n269), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT95), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n509), .A2(new_n512), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n356), .A2(new_n361), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n294), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n566), .A2(new_n555), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n284), .A2(new_n570), .A3(new_n285), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n281), .A2(KEYINPUT96), .A3(new_n283), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n289), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n442), .A2(KEYINPUT33), .A3(new_n443), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n453), .B2(new_n441), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n575), .A2(new_n577), .A3(G478), .A4(new_n269), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n269), .B1(new_n453), .B2(new_n441), .ZN(new_n579));
  NAND2_X1  g393(.A1(KEYINPUT97), .A2(G478), .ZN(new_n580));
  OR2_X1    g394(.A1(KEYINPUT97), .A2(G478), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT98), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n578), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n416), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n463), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n574), .A2(new_n589), .A3(KEYINPUT99), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n571), .A2(new_n590), .A3(new_n289), .A4(new_n572), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(new_n588), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n569), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  NAND3_X1  g412(.A1(new_n407), .A2(KEYINPUT100), .A3(new_n410), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n410), .A2(KEYINPUT100), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n415), .ZN(new_n601));
  INV_X1    g415(.A(new_n456), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n593), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n569), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n538), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n553), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n549), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n565), .B(new_n610), .C1(new_n561), .C2(new_n563), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT101), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n465), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT37), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n525), .ZN(G12));
  NAND2_X1  g429(.A1(new_n518), .A2(new_n519), .ZN(new_n616));
  INV_X1    g430(.A(new_n502), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n458), .B1(new_n462), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n599), .A2(new_n600), .A3(new_n415), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n549), .A2(new_n609), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n622), .A2(new_n623), .A3(new_n602), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n618), .A2(new_n624), .A3(new_n362), .A4(new_n574), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XNOR2_X1  g440(.A(new_n288), .B(KEYINPUT38), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n485), .B1(new_n487), .B2(new_n493), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n628), .A2(G902), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n479), .A2(new_n485), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n616), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n416), .A2(new_n456), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n627), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n610), .A2(new_n290), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n620), .B(KEYINPUT39), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n362), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT40), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n637), .A2(KEYINPUT40), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n634), .A2(new_n635), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n210), .ZN(G45));
  NAND4_X1  g455(.A1(new_n610), .A2(new_n416), .A3(new_n587), .A4(new_n621), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n618), .A2(new_n362), .A3(new_n643), .A4(new_n574), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  NAND2_X1  g459(.A1(new_n354), .A2(new_n269), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G469), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n356), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n649), .A3(G469), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n295), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n595), .A2(new_n651), .A3(new_n556), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT103), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n595), .A2(new_n651), .A3(new_n654), .A4(new_n556), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G113), .ZN(G15));
  NAND3_X1  g472(.A1(new_n651), .A2(new_n556), .A3(new_n603), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G116), .ZN(G18));
  INV_X1    g474(.A(new_n464), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n520), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n651), .A2(new_n662), .A3(new_n574), .A4(new_n610), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  NOR2_X1   g478(.A1(new_n593), .A2(new_n602), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT104), .B(G472), .Z(new_n666));
  NOR2_X1   g480(.A1(new_n559), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n497), .A2(new_n500), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n485), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n511), .B1(new_n669), .B2(new_n507), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n667), .A2(new_n670), .A3(new_n555), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n651), .A2(new_n416), .A3(new_n665), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  NOR3_X1   g487(.A1(new_n642), .A2(new_n670), .A3(new_n667), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n651), .A2(new_n574), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(G125), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G27));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n588), .A2(new_n620), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n568), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n288), .A2(new_n289), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n362), .A2(KEYINPUT106), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT107), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n688), .A3(new_n684), .A4(new_n685), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n678), .B(new_n680), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n555), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n513), .A2(new_n516), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n691), .B1(new_n502), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT106), .B1(new_n567), .B2(new_n294), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n681), .B(new_n295), .C1(new_n356), .C2(new_n361), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n688), .B1(new_n697), .B2(new_n684), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT107), .A4(new_n683), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n556), .B(new_n679), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n690), .A2(new_n694), .B1(new_n678), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G131), .ZN(G33));
  INV_X1    g517(.A(new_n556), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n687), .B2(new_n689), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n622), .A2(new_n602), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G134), .ZN(G36));
  NAND3_X1  g522(.A1(new_n587), .A2(new_n411), .A3(new_n415), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT111), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT43), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(KEYINPUT44), .A3(new_n566), .A4(new_n610), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n360), .B2(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT109), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n360), .A2(KEYINPUT45), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n717), .B(G469), .C1(new_n360), .C2(KEYINPUT45), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(G469), .A2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n719), .A2(new_n725), .A3(KEYINPUT46), .A4(new_n720), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n724), .A3(new_n356), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n294), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n711), .A2(new_n566), .A3(new_n610), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n729), .A3(new_n636), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n728), .B1(new_n735), .B2(KEYINPUT47), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(KEYINPUT47), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n735), .A2(KEYINPUT47), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n727), .B(new_n294), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n684), .A2(new_n555), .A3(new_n520), .A4(new_n679), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT113), .Z(new_n741));
  NAND3_X1  g555(.A1(new_n736), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  AOI21_X1  g557(.A(new_n610), .B1(new_n616), .B2(new_n631), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n573), .A2(new_n633), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n362), .A3(new_n621), .A4(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n675), .A2(new_n746), .A3(new_n625), .A4(new_n644), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n625), .A2(new_n644), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(KEYINPUT52), .A3(new_n675), .A4(new_n746), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n557), .A2(new_n613), .A3(new_n659), .A4(new_n672), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n456), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT115), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n411), .A3(new_n415), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n588), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n291), .A2(new_n759), .A3(new_n590), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n568), .A2(new_n555), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n565), .A4(new_n564), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n663), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n653), .B2(new_n655), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n752), .A2(new_n753), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n701), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n674), .B1(new_n698), .B2(new_n699), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n687), .A2(new_n689), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT116), .A3(new_n674), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n568), .A2(new_n520), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n623), .A2(new_n757), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n683), .A2(new_n622), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n705), .B2(new_n706), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n773), .B1(new_n772), .B2(new_n779), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n766), .B(KEYINPUT53), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT116), .B1(new_n770), .B2(new_n674), .ZN(new_n784));
  INV_X1    g598(.A(new_n674), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n768), .B(new_n785), .C1(new_n687), .C2(new_n689), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n707), .A2(new_n777), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT117), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n791), .B2(new_n766), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n651), .A2(new_n684), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT119), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n711), .A2(new_n458), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n797), .A2(new_n623), .A3(new_n670), .A4(new_n667), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n632), .A2(new_n458), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n691), .A3(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n416), .A3(new_n587), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n651), .A2(new_n671), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n290), .A3(new_n627), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT50), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n798), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n796), .A2(new_n671), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n684), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n648), .A2(new_n650), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT114), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n809), .A2(new_n294), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n736), .A2(new_n739), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT118), .B1(new_n736), .B2(new_n739), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n807), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n805), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n810), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n807), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n816), .A2(new_n817), .B1(new_n805), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n766), .B1(new_n780), .B2(new_n781), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n782), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n793), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n806), .A2(new_n574), .A3(new_n651), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n795), .A2(new_n691), .A3(new_n589), .A4(new_n799), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n457), .A2(G953), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT48), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n797), .B2(new_n693), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n795), .A2(new_n796), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(KEYINPUT48), .A3(new_n694), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT120), .A4(new_n829), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n834), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT121), .Z(new_n839));
  OAI22_X1  g653(.A1(new_n826), .A2(new_n839), .B1(G952), .B2(G953), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n809), .B(KEYINPUT49), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n709), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n555), .A2(new_n295), .A3(new_n290), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n632), .A3(new_n627), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(G75));
  NAND2_X1  g659(.A1(new_n457), .A2(G953), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT122), .Z(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n269), .B1(new_n823), .B2(new_n782), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n849), .B2(G210), .ZN(new_n850));
  INV_X1    g664(.A(new_n264), .ZN(new_n851));
  INV_X1    g665(.A(new_n265), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n267), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n224), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT55), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(G210), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n858), .B(new_n269), .C1(new_n823), .C2(new_n782), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n855), .B1(new_n859), .B2(KEYINPUT56), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n848), .B1(new_n857), .B2(new_n860), .ZN(G51));
  XOR2_X1   g675(.A(new_n720), .B(KEYINPUT57), .Z(new_n862));
  AND3_X1   g676(.A1(new_n823), .A2(new_n824), .A3(new_n782), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n824), .B1(new_n823), .B2(new_n782), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n354), .ZN(new_n866));
  INV_X1    g680(.A(new_n719), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n848), .B1(new_n866), .B2(new_n868), .ZN(G54));
  NAND3_X1  g683(.A1(new_n849), .A2(KEYINPUT58), .A3(G475), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n404), .ZN(new_n871));
  INV_X1    g685(.A(new_n404), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n849), .A2(KEYINPUT58), .A3(G475), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n848), .B1(new_n871), .B2(new_n873), .ZN(G60));
  NAND2_X1  g688(.A1(G478), .A2(G902), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT59), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n863), .B2(new_n864), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n575), .A2(new_n577), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n878), .B(new_n876), .C1(new_n863), .C2(new_n864), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n848), .B1(new_n880), .B2(new_n881), .ZN(G63));
  NAND2_X1  g696(.A1(G217), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT60), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n783), .B2(new_n792), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n848), .B1(new_n886), .B2(new_n550), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n608), .B(new_n885), .C1(new_n783), .C2(new_n792), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(KEYINPUT123), .C2(KEYINPUT61), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n884), .B1(new_n823), .B2(new_n782), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n888), .B(new_n847), .C1(new_n551), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT61), .B1(new_n888), .B2(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(G66));
  NAND2_X1  g708(.A1(new_n753), .A2(new_n764), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(G953), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n218), .B1(new_n460), .B2(new_n219), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(KEYINPUT124), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n853), .B1(G898), .B2(new_n218), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(G69));
  NAND2_X1  g716(.A1(new_n491), .A2(new_n492), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n377), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT125), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n750), .A2(new_n675), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n640), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT62), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n733), .A2(new_n742), .ZN(new_n909));
  INV_X1    g723(.A(new_n637), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n556), .A3(new_n684), .A4(new_n759), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT126), .Z(new_n912));
  NOR3_X1   g726(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n905), .B1(new_n913), .B2(G953), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n619), .A2(new_n218), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n733), .A2(new_n742), .A3(new_n707), .ZN(new_n916));
  INV_X1    g730(.A(new_n701), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n729), .A2(new_n636), .A3(new_n694), .A4(new_n745), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n906), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n904), .B1(new_n919), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G72));
  NAND2_X1  g737(.A1(G472), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT63), .Z(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n919), .B2(new_n895), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n494), .A2(new_n498), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT127), .B(new_n925), .C1(new_n919), .C2(new_n895), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n913), .A2(new_n896), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n925), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n628), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n847), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n925), .B1(new_n494), .B2(new_n498), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n628), .B(new_n936), .C1(new_n823), .C2(new_n782), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(G57));
endmodule


