

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U321 ( .A(n307), .B(n306), .Z(n525) );
  XOR2_X1 U322 ( .A(KEYINPUT28), .B(n474), .Z(n527) );
  XOR2_X1 U323 ( .A(n350), .B(n401), .Z(n289) );
  XOR2_X1 U324 ( .A(G43GAT), .B(G99GAT), .Z(n290) );
  XNOR2_X1 U325 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U326 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U327 ( .A(n308), .B(n290), .ZN(n304) );
  XNOR2_X1 U328 ( .A(n414), .B(n413), .ZN(n566) );
  XNOR2_X1 U329 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U330 ( .A(KEYINPUT119), .B(n477), .ZN(n563) );
  INV_X1 U331 ( .A(G43GAT), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n496) );
  XNOR2_X1 U333 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n478) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U335 ( .A(n479), .B(n478), .ZN(G1350GAT) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U337 ( .A(G176GAT), .B(KEYINPUT84), .Z(n292) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n307) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G127GAT), .Z(n350) );
  INV_X1 U341 ( .A(KEYINPUT19), .ZN(n293) );
  NAND2_X1 U342 ( .A1(KEYINPUT18), .A2(n293), .ZN(n296) );
  INV_X1 U343 ( .A(KEYINPUT18), .ZN(n294) );
  NAND2_X1 U344 ( .A1(n294), .A2(KEYINPUT19), .ZN(n295) );
  NAND2_X1 U345 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n401) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n289), .B(n299), .ZN(n301) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n300), .B(KEYINPUT0), .ZN(n370) );
  XOR2_X1 U352 ( .A(n301), .B(n370), .Z(n303) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(KEYINPUT65), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n308) );
  XOR2_X1 U356 ( .A(G57GAT), .B(KEYINPUT13), .Z(n343) );
  XNOR2_X1 U357 ( .A(n308), .B(n343), .ZN(n323) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n309), .B(KEYINPUT73), .ZN(n424) );
  XOR2_X1 U360 ( .A(n424), .B(KEYINPUT33), .Z(n311) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n321) );
  XOR2_X1 U367 ( .A(G78GAT), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n398) );
  XOR2_X1 U370 ( .A(G64GAT), .B(G92GAT), .Z(n319) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n405) );
  XNOR2_X1 U373 ( .A(n398), .B(n405), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n574) );
  XOR2_X1 U376 ( .A(G197GAT), .B(G22GAT), .Z(n325) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(G141GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n327) );
  XNOR2_X1 U380 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n341) );
  XOR2_X1 U383 ( .A(G1GAT), .B(KEYINPUT70), .Z(n351) );
  XOR2_X1 U384 ( .A(G113GAT), .B(G15GAT), .Z(n331) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G50GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U387 ( .A(n351), .B(n332), .Z(n334) );
  NAND2_X1 U388 ( .A1(G229GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n335), .B(KEYINPUT30), .Z(n339) );
  XOR2_X1 U391 ( .A(G29GAT), .B(G43GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n434) );
  XNOR2_X1 U394 ( .A(n434), .B(KEYINPUT69), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U396 ( .A(n341), .B(n340), .Z(n568) );
  INV_X1 U397 ( .A(n568), .ZN(n554) );
  NAND2_X1 U398 ( .A1(n574), .A2(n554), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(KEYINPUT76), .ZN(n483) );
  XOR2_X1 U400 ( .A(G8GAT), .B(G183GAT), .Z(n404) );
  XOR2_X1 U401 ( .A(n404), .B(n343), .Z(n345) );
  XNOR2_X1 U402 ( .A(G71GAT), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  XOR2_X1 U405 ( .A(n385), .B(KEYINPUT82), .Z(n347) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U408 ( .A(n349), .B(n348), .Z(n353) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n361) );
  XOR2_X1 U411 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n355) );
  XNOR2_X1 U412 ( .A(G78GAT), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U414 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n357) );
  XNOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U417 ( .A(n359), .B(n358), .Z(n360) );
  XOR2_X1 U418 ( .A(n361), .B(n360), .Z(n579) );
  XOR2_X1 U419 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n363) );
  XNOR2_X1 U420 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(G155GAT), .Z(n365) );
  XNOR2_X1 U423 ( .A(G120GAT), .B(G148GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n382) );
  XOR2_X1 U426 ( .A(G85GAT), .B(G162GAT), .Z(n369) );
  XNOR2_X1 U427 ( .A(G29GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U429 ( .A(n370), .B(G57GAT), .Z(n372) );
  NAND2_X1 U430 ( .A1(G225GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n380) );
  XNOR2_X1 U433 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(KEYINPUT2), .ZN(n393) );
  XOR2_X1 U435 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n377) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n393), .B(n378), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n473) );
  XOR2_X1 U441 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n384) );
  XNOR2_X1 U442 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n387) );
  XOR2_X1 U445 ( .A(G50GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U446 ( .A(n433), .B(n385), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U448 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U451 ( .A(n392), .B(KEYINPUT22), .Z(n395) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT23), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U454 ( .A(G211GAT), .B(KEYINPUT21), .Z(n397) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(G218GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n406) );
  XOR2_X1 U457 ( .A(n406), .B(n398), .Z(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n474) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(n401), .Z(n403) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n410) );
  XOR2_X1 U462 ( .A(n405), .B(n404), .Z(n408) );
  XOR2_X1 U463 ( .A(G36GAT), .B(G190GAT), .Z(n430) );
  XNOR2_X1 U464 ( .A(n406), .B(n430), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n515) );
  NAND2_X1 U467 ( .A1(n525), .A2(n515), .ZN(n411) );
  NAND2_X1 U468 ( .A1(n474), .A2(n411), .ZN(n412) );
  XOR2_X1 U469 ( .A(KEYINPUT25), .B(n412), .Z(n416) );
  NOR2_X1 U470 ( .A1(n525), .A2(n474), .ZN(n414) );
  XNOR2_X1 U471 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n515), .B(KEYINPUT27), .ZN(n418) );
  NAND2_X1 U473 ( .A1(n566), .A2(n418), .ZN(n415) );
  NAND2_X1 U474 ( .A1(n416), .A2(n415), .ZN(n417) );
  NAND2_X1 U475 ( .A1(n473), .A2(n417), .ZN(n422) );
  INV_X1 U476 ( .A(n527), .ZN(n420) );
  INV_X1 U477 ( .A(n473), .ZN(n513) );
  NAND2_X1 U478 ( .A1(n513), .A2(n418), .ZN(n522) );
  NOR2_X1 U479 ( .A1(n525), .A2(n522), .ZN(n419) );
  NAND2_X1 U480 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND2_X1 U481 ( .A1(n422), .A2(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(KEYINPUT95), .B(n423), .Z(n481) );
  NAND2_X1 U483 ( .A1(n579), .A2(n481), .ZN(n450) );
  NAND2_X1 U484 ( .A1(n424), .A2(KEYINPUT10), .ZN(n428) );
  INV_X1 U485 ( .A(n424), .ZN(n426) );
  INV_X1 U486 ( .A(KEYINPUT10), .ZN(n425) );
  NAND2_X1 U487 ( .A1(n426), .A2(n425), .ZN(n427) );
  NAND2_X1 U488 ( .A1(n428), .A2(n427), .ZN(n432) );
  AND2_X1 U489 ( .A1(G232GAT), .A2(G233GAT), .ZN(n429) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U492 ( .A(G92GAT), .B(KEYINPUT67), .Z(n438) );
  XNOR2_X1 U493 ( .A(G134GAT), .B(G218GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n448) );
  XOR2_X1 U496 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n442) );
  XNOR2_X1 U497 ( .A(G106GAT), .B(KEYINPUT66), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U499 ( .A(KEYINPUT78), .B(KEYINPUT64), .Z(n444) );
  XNOR2_X1 U500 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X2 U503 ( .A(n448), .B(n447), .ZN(n562) );
  XOR2_X1 U504 ( .A(n562), .B(KEYINPUT98), .Z(n449) );
  XNOR2_X1 U505 ( .A(n449), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U506 ( .A1(n450), .A2(n583), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(KEYINPUT37), .ZN(n512) );
  NOR2_X1 U508 ( .A1(n483), .A2(n512), .ZN(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT99), .B(KEYINPUT38), .Z(n452) );
  NAND2_X1 U510 ( .A1(n525), .A2(n496), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n455) );
  INV_X1 U512 ( .A(n579), .ZN(n549) );
  XNOR2_X1 U513 ( .A(KEYINPUT41), .B(n574), .ZN(n544) );
  NAND2_X1 U514 ( .A1(n554), .A2(n544), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT46), .B(n458), .ZN(n460) );
  INV_X1 U516 ( .A(n562), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n549), .A2(n461), .ZN(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT47), .B(n462), .Z(n468) );
  NOR2_X1 U520 ( .A1(n579), .A2(n583), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT45), .B(n463), .ZN(n465) );
  AND2_X1 U522 ( .A1(n574), .A2(n568), .ZN(n464) );
  AND2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(KEYINPUT108), .B(n466), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT48), .B(n469), .ZN(n523) );
  XOR2_X1 U527 ( .A(n515), .B(KEYINPUT118), .Z(n470) );
  NOR2_X1 U528 ( .A1(n523), .A2(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT54), .B(n471), .ZN(n472) );
  AND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n567) );
  NAND2_X1 U531 ( .A1(n567), .A2(n474), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT55), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n476), .A2(n525), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n549), .A2(n563), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n485) );
  NOR2_X1 U536 ( .A1(n579), .A2(n562), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n480), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n500) );
  NOR2_X1 U539 ( .A1(n483), .A2(n500), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n491), .A2(n513), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n486), .Z(G1324GAT) );
  XOR2_X1 U543 ( .A(G8GAT), .B(KEYINPUT97), .Z(n488) );
  NAND2_X1 U544 ( .A1(n491), .A2(n515), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U547 ( .A1(n491), .A2(n525), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n527), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U552 ( .A1(n513), .A2(n496), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n515), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n498) );
  NAND2_X1 U557 ( .A1(n496), .A2(n527), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(n544), .Z(n557) );
  NAND2_X1 U562 ( .A1(n568), .A2(n557), .ZN(n511) );
  NOR2_X1 U563 ( .A1(n511), .A2(n500), .ZN(n507) );
  NAND2_X1 U564 ( .A1(n513), .A2(n507), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n515), .A2(n507), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U570 ( .A1(n507), .A2(n525), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U573 ( .A1(n507), .A2(n527), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n513), .A2(n518), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n518), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n525), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n527), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U588 ( .A(KEYINPUT109), .B(n524), .Z(n540) );
  NAND2_X1 U589 ( .A1(n525), .A2(n540), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n536), .A2(n554), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n531) );
  NAND2_X1 U595 ( .A1(n536), .A2(n557), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT111), .Z(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n549), .A2(n536), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT51), .B(KEYINPUT113), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n562), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  XOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U607 ( .A1(n540), .A2(n566), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n541), .Z(n552) );
  NAND2_X1 U609 ( .A1(n554), .A2(n552), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n548) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U613 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n562), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n563), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n582) );
  NOR2_X1 U633 ( .A1(n568), .A2(n582), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT123), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n582), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

