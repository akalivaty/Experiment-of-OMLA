

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586;

  XOR2_X1 U327 ( .A(G204GAT), .B(G78GAT), .Z(n295) );
  INV_X1 U328 ( .A(KEYINPUT47), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n445), .B(n295), .ZN(n380) );
  XNOR2_X1 U330 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U331 ( .A(n422), .B(n478), .ZN(n550) );
  XNOR2_X1 U332 ( .A(n456), .B(G176GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U337 ( .A(n298), .B(G99GAT), .Z(n300) );
  XOR2_X1 U338 ( .A(G134GAT), .B(KEYINPUT0), .Z(n448) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(n448), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n306) );
  XOR2_X1 U341 ( .A(KEYINPUT17), .B(KEYINPUT84), .Z(n302) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n341) );
  XOR2_X1 U344 ( .A(n341), .B(KEYINPUT82), .Z(n304) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U347 ( .A(n306), .B(n305), .Z(n314) );
  XOR2_X1 U348 ( .A(G183GAT), .B(G15GAT), .Z(n308) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(G113GAT), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U351 ( .A(G71GAT), .B(G127GAT), .Z(n310) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(G176GAT), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U354 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U355 ( .A(n314), .B(n313), .ZN(n532) );
  XOR2_X1 U356 ( .A(KEYINPUT88), .B(G218GAT), .Z(n316) );
  XNOR2_X1 U357 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U358 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U359 ( .A(KEYINPUT87), .B(n317), .Z(n349) );
  XOR2_X1 U360 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n319) );
  XNOR2_X1 U361 ( .A(G162GAT), .B(KEYINPUT89), .ZN(n318) );
  XNOR2_X1 U362 ( .A(n319), .B(n318), .ZN(n447) );
  XOR2_X1 U363 ( .A(G155GAT), .B(G78GAT), .Z(n383) );
  XOR2_X1 U364 ( .A(n447), .B(n383), .Z(n321) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U367 ( .A(n349), .B(n322), .ZN(n335) );
  XOR2_X1 U368 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n324) );
  XNOR2_X1 U369 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U371 ( .A(G148GAT), .B(KEYINPUT90), .Z(n326) );
  XNOR2_X1 U372 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U374 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U375 ( .A(G22GAT), .B(G197GAT), .Z(n330) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U380 ( .A(n335), .B(n334), .ZN(n470) );
  XOR2_X1 U381 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n337) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U383 ( .A(n337), .B(n336), .ZN(n340) );
  XOR2_X1 U384 ( .A(G64GAT), .B(KEYINPUT78), .Z(n339) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G92GAT), .ZN(n338) );
  XNOR2_X1 U386 ( .A(n339), .B(n338), .ZN(n377) );
  XOR2_X1 U387 ( .A(n340), .B(n377), .Z(n343) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U389 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U390 ( .A(G183GAT), .B(G211GAT), .Z(n395) );
  XOR2_X1 U391 ( .A(n344), .B(n395), .Z(n347) );
  XNOR2_X1 U392 ( .A(G169GAT), .B(G197GAT), .ZN(n345) );
  XNOR2_X1 U393 ( .A(n345), .B(G8GAT), .ZN(n367) );
  XOR2_X1 U394 ( .A(G190GAT), .B(KEYINPUT80), .Z(n398) );
  XNOR2_X1 U395 ( .A(n367), .B(n398), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U397 ( .A(n349), .B(n348), .ZN(n519) );
  INV_X1 U398 ( .A(KEYINPUT117), .ZN(n421) );
  XOR2_X1 U399 ( .A(G43GAT), .B(G29GAT), .Z(n351) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U402 ( .A(n352), .B(KEYINPUT73), .Z(n354) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n412) );
  XOR2_X1 U405 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n356) );
  XNOR2_X1 U406 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U408 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n358) );
  XNOR2_X1 U409 ( .A(KEYINPUT74), .B(KEYINPUT68), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U411 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U412 ( .A(KEYINPUT29), .B(KEYINPUT72), .Z(n362) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U415 ( .A(KEYINPUT30), .B(n363), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G22GAT), .Z(n388) );
  XOR2_X1 U418 ( .A(n366), .B(n388), .Z(n369) );
  XOR2_X1 U419 ( .A(G113GAT), .B(G141GAT), .Z(n436) );
  XNOR2_X1 U420 ( .A(n436), .B(n367), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U422 ( .A(n412), .B(n370), .Z(n570) );
  XNOR2_X1 U423 ( .A(n570), .B(KEYINPUT76), .ZN(n558) );
  INV_X1 U424 ( .A(KEYINPUT116), .ZN(n418) );
  XOR2_X1 U425 ( .A(KEYINPUT77), .B(KEYINPUT13), .Z(n372) );
  XNOR2_X1 U426 ( .A(G71GAT), .B(G57GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U428 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n374) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U431 ( .A(n375), .B(KEYINPUT32), .Z(n379) );
  XNOR2_X1 U432 ( .A(G99GAT), .B(G106GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n376), .B(G85GAT), .ZN(n399) );
  XNOR2_X1 U434 ( .A(n377), .B(n399), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U436 ( .A(G120GAT), .B(G148GAT), .Z(n445) );
  XOR2_X1 U437 ( .A(n384), .B(n382), .Z(n575) );
  XOR2_X1 U438 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n415) );
  XOR2_X1 U439 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n387), .B(G64GAT), .ZN(n390) );
  XOR2_X1 U443 ( .A(G8GAT), .B(n388), .Z(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n394) );
  XOR2_X1 U445 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n392) );
  XNOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n397) );
  XOR2_X1 U449 ( .A(G1GAT), .B(G127GAT), .Z(n435) );
  XNOR2_X1 U450 ( .A(n435), .B(n395), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n579) );
  XNOR2_X1 U452 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n413) );
  XOR2_X1 U453 ( .A(n399), .B(n398), .Z(n401) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(G162GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n403) );
  NAND2_X1 U457 ( .A1(G232GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U460 ( .A(KEYINPUT79), .B(KEYINPUT66), .Z(n407) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n408), .B(KEYINPUT9), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n459) );
  XNOR2_X1 U466 ( .A(n413), .B(n459), .ZN(n581) );
  NAND2_X1 U467 ( .A1(n579), .A2(n581), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  NOR2_X1 U469 ( .A1(n575), .A2(n416), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n419) );
  NOR2_X1 U471 ( .A1(n558), .A2(n419), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n429) );
  INV_X1 U473 ( .A(n459), .ZN(n564) );
  XNOR2_X1 U474 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n422) );
  INV_X1 U475 ( .A(n575), .ZN(n478) );
  NAND2_X1 U476 ( .A1(n570), .A2(n550), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n423), .B(KEYINPUT46), .ZN(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT115), .B(n579), .ZN(n562) );
  NAND2_X1 U479 ( .A1(n424), .A2(n562), .ZN(n425) );
  NOR2_X1 U480 ( .A1(n564), .A2(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  NOR2_X1 U482 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U483 ( .A(KEYINPUT48), .B(n430), .ZN(n530) );
  NOR2_X1 U484 ( .A1(n519), .A2(n530), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT54), .ZN(n453) );
  XOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n433) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(KEYINPUT1), .B(n434), .ZN(n452) );
  XOR2_X1 U490 ( .A(KEYINPUT92), .B(n435), .Z(n438) );
  XNOR2_X1 U491 ( .A(n436), .B(G155GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U493 ( .A(n439), .B(G85GAT), .Z(n444) );
  XOR2_X1 U494 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n441) );
  XNOR2_X1 U495 ( .A(G57GAT), .B(KEYINPUT93), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n469) );
  XNOR2_X1 U503 ( .A(KEYINPUT95), .B(n469), .ZN(n517) );
  NAND2_X1 U504 ( .A1(n453), .A2(n517), .ZN(n569) );
  NOR2_X1 U505 ( .A1(n470), .A2(n569), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NOR2_X2 U507 ( .A1(n532), .A2(n455), .ZN(n565) );
  NAND2_X1 U508 ( .A1(n565), .A2(n550), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  NAND2_X1 U510 ( .A1(n579), .A2(n459), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n460), .ZN(n476) );
  NOR2_X1 U512 ( .A1(n532), .A2(n519), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n470), .A2(n461), .ZN(n462) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n462), .Z(n467) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(n519), .ZN(n471) );
  NAND2_X1 U517 ( .A1(n470), .A2(n532), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT26), .ZN(n465) );
  XNOR2_X1 U519 ( .A(KEYINPUT100), .B(n465), .ZN(n568) );
  NOR2_X1 U520 ( .A1(n471), .A2(n568), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n469), .A2(n468), .ZN(n475) );
  XOR2_X1 U523 ( .A(n470), .B(KEYINPUT28), .Z(n531) );
  NAND2_X1 U524 ( .A1(n532), .A2(n531), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n471), .A2(n517), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT99), .ZN(n529) );
  NOR2_X1 U527 ( .A1(n473), .A2(n529), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n487) );
  NOR2_X1 U529 ( .A1(n476), .A2(n487), .ZN(n477) );
  XNOR2_X1 U530 ( .A(n477), .B(KEYINPUT101), .ZN(n503) );
  NAND2_X1 U531 ( .A1(n558), .A2(n478), .ZN(n490) );
  NOR2_X1 U532 ( .A1(n503), .A2(n490), .ZN(n479) );
  XOR2_X1 U533 ( .A(KEYINPUT102), .B(n479), .Z(n485) );
  NOR2_X1 U534 ( .A1(n485), .A2(n517), .ZN(n480) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(n480), .Z(n481) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n485), .A2(n519), .ZN(n482) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n484) );
  NOR2_X1 U540 ( .A1(n532), .A2(n485), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n531), .A2(n485), .ZN(n486) );
  XOR2_X1 U543 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  NOR2_X1 U544 ( .A1(n579), .A2(n487), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n581), .A2(n488), .ZN(n489) );
  XOR2_X1 U546 ( .A(KEYINPUT37), .B(n489), .Z(n514) );
  NOR2_X1 U547 ( .A1(n490), .A2(n514), .ZN(n491) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n491), .Z(n497) );
  NOR2_X1 U549 ( .A1(n497), .A2(n517), .ZN(n493) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n497), .A2(n519), .ZN(n494) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n532), .A2(n497), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(n495), .Z(n496) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n531), .A2(n497), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  INV_X1 U561 ( .A(n570), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n550), .A2(n501), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT106), .ZN(n515) );
  OR2_X1 U564 ( .A1(n515), .A2(n503), .ZN(n510) );
  NOR2_X1 U565 ( .A1(n517), .A2(n510), .ZN(n505) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n510), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n532), .A2(n510), .ZN(n509) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n531), .A2(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  NOR2_X1 U578 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT110), .B(n516), .Z(n525) );
  NOR2_X1 U580 ( .A1(n525), .A2(n517), .ZN(n518) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n525), .A2(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n532), .A2(n525), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n546), .A2(n531), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT118), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n558), .A2(n542), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U600 ( .A1(n542), .A2(n550), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  INV_X1 U603 ( .A(n542), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n539), .A2(n562), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U608 ( .A1(n564), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT121), .Z(n549) );
  INV_X1 U612 ( .A(n546), .ZN(n547) );
  NOR2_X1 U613 ( .A1(n568), .A2(n547), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n555), .A2(n570), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n555), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n579), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n564), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT122), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  XOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT123), .Z(n560) );
  NAND2_X1 U626 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  INV_X1 U628 ( .A(n565), .ZN(n561) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .Z(n572) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n582), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n586) );
  XOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n584) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1355GAT) );
endmodule

