//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n466), .B1(new_n461), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n468), .B1(new_n462), .B2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n480), .B(new_n484), .C1(G136), .C2(new_n464), .ZN(G162));
  NAND3_X1  g060(.A1(new_n473), .A2(G138), .A3(new_n468), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n488), .A2(new_n489), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT71), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT71), .A2(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n501), .A2(new_n506), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n501), .A2(G543), .A3(new_n509), .A4(new_n511), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n498), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n517), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n506), .A2(G62), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n506), .A2(new_n523), .A3(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n500), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT71), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT75), .B1(new_n525), .B2(new_n529), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n518), .A2(new_n520), .B1(new_n532), .B2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n516), .A2(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n513), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  INV_X1    g115(.A(new_n505), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n504), .A2(KEYINPUT76), .A3(new_n505), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(G63), .A3(G651), .ZN(new_n546));
  AND4_X1   g121(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n546), .ZN(G168));
  AND2_X1   g122(.A1(new_n511), .A2(new_n509), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n548), .A2(G52), .A3(G543), .A4(new_n501), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n548), .A2(G90), .A3(new_n506), .A4(new_n501), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n543), .A2(new_n544), .A3(G64), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n528), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT77), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n549), .A2(new_n550), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n554), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n561), .A2(new_n515), .B1(new_n512), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n543), .A2(new_n544), .A3(G56), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n528), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NOR3_X1   g147(.A1(new_n526), .A2(new_n527), .A3(new_n508), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n511), .A2(new_n509), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n515), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G91), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n512), .A2(new_n581), .B1(new_n582), .B2(new_n510), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  NAND4_X1  g161(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n546), .ZN(G286));
  NAND2_X1  g162(.A1(new_n513), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n545), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n516), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI21_X1  g166(.A(KEYINPUT78), .B1(new_n506), .B2(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G73), .B2(G543), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n506), .A2(KEYINPUT78), .A3(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n528), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n515), .B1(new_n512), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n545), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n528), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n604), .A2(new_n515), .B1(new_n512), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND4_X1  g183(.A1(new_n575), .A2(KEYINPUT10), .A3(G92), .A4(new_n506), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n515), .A2(new_n614), .B1(new_n615), .B2(new_n510), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g195(.A(new_n619), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n583), .B1(new_n579), .B2(new_n577), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(G297));
  XOR2_X1   g199(.A(G297), .B(KEYINPUT80), .Z(G280));
  AOI21_X1  g200(.A(new_n616), .B1(new_n612), .B2(new_n609), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  OAI21_X1  g203(.A(KEYINPUT82), .B1(new_n567), .B2(G868), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n618), .B2(G559), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(KEYINPUT81), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  MUX2_X1   g209(.A(KEYINPUT82), .B(new_n629), .S(new_n634), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n470), .A2(new_n473), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n464), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n481), .A2(G123), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  OAI211_X1 g223(.A(new_n642), .B(new_n648), .C1(G2100), .C2(new_n640), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n672), .B(new_n669), .C1(new_n665), .C2(new_n667), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n665), .A3(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n683), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n684), .B1(new_n681), .B2(new_n685), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  XOR2_X1   g272(.A(KEYINPUT87), .B(G29), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G35), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G162), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT29), .Z(new_n702));
  INV_X1    g277(.A(G2090), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G4), .A2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n618), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT91), .B(G1348), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n698), .A2(G26), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  OAI211_X1 g287(.A(G140), .B(new_n468), .C1(new_n490), .C2(new_n491), .ZN(new_n713));
  OAI211_X1 g288(.A(G128), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(G116), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G2105), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n717), .A3(G2104), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n714), .A3(new_n721), .A4(new_n718), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n712), .B1(G29), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2067), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n704), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  OAI22_X1  g301(.A1(new_n702), .A2(new_n703), .B1(new_n709), .B2(new_n708), .ZN(new_n727));
  NOR3_X1   g302(.A1(KEYINPUT94), .A2(G5), .A3(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT94), .B1(G5), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n728), .B(new_n730), .C1(G171), .C2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT95), .B(G1961), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n699), .A2(G27), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n699), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2078), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n567), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT92), .B(G1341), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n737), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G20), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT23), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n733), .A2(new_n734), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(G34), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n698), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  INV_X1    g330(.A(G32), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n470), .A2(G105), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n473), .A2(G141), .A3(new_n468), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n473), .A2(G129), .A3(G2105), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT26), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n754), .A2(new_n755), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  INV_X1    g345(.A(G33), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n473), .A2(G139), .A3(new_n468), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n774));
  NAND2_X1  g349(.A1(G103), .A2(G2104), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n473), .A2(G127), .ZN(new_n781));
  NAND2_X1  g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2105), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n772), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G2072), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n754), .A2(new_n755), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT30), .A2(G28), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT30), .A2(G28), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(G29), .B2(new_n792), .C1(new_n647), .C2(new_n698), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n770), .A2(new_n787), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n707), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n707), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1966), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n726), .A2(new_n727), .A3(new_n748), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  NOR2_X1   g375(.A1(G303), .A2(new_n707), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G22), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n801), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n707), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n707), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n804), .A2(new_n805), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G6), .A2(G16), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n599), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  INV_X1    g389(.A(G1981), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n811), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n699), .A2(G25), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n473), .A2(G131), .A3(new_n468), .ZN(new_n822));
  OAI211_X1 g397(.A(G119), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(new_n699), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n828), .B(new_n829), .Z(new_n830));
  AOI21_X1  g405(.A(new_n707), .B1(G290), .B2(KEYINPUT88), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(KEYINPUT88), .B2(G290), .ZN(new_n832));
  INV_X1    g407(.A(G24), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(G16), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n830), .B1(new_n834), .B2(G1986), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G1986), .B2(new_n834), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n818), .A2(new_n820), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT89), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(KEYINPUT89), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n800), .B1(new_n840), .B2(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  NAND3_X1  g418(.A1(new_n543), .A2(new_n544), .A3(G67), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n529), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(KEYINPUT97), .A3(new_n529), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n566), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n516), .A2(G43), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n513), .A2(G81), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(KEYINPUT98), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n563), .B2(new_n566), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n512), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n515), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n851), .A2(new_n855), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT97), .B1(new_n846), .B2(new_n529), .ZN(new_n864));
  AOI211_X1 g439(.A(new_n848), .B(new_n528), .C1(new_n844), .C2(new_n845), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n567), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n856), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT38), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n626), .A2(G559), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n866), .A2(G860), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n877), .ZN(G145));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n766), .A2(new_n780), .A3(new_n784), .ZN(new_n880));
  AOI22_X1  g455(.A1(G141), .A2(new_n464), .B1(new_n470), .B2(G105), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n481), .A2(G129), .B1(new_n763), .B2(new_n764), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n468), .B1(new_n781), .B2(new_n782), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n779), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n723), .A2(new_n496), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT4), .B1(new_n464), .B2(G138), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n492), .A2(new_n495), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n489), .A2(new_n889), .B1(new_n720), .B2(new_n722), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n885), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n723), .A2(new_n496), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n889), .A2(new_n720), .A3(new_n489), .A4(new_n722), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n884), .A4(new_n880), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n637), .B(new_n638), .Z(new_n897));
  OAI211_X1 g472(.A(G130), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT99), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n473), .A2(new_n900), .A3(G130), .A4(G2105), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n903));
  INV_X1    g478(.A(G118), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n903), .A2(KEYINPUT100), .B1(new_n904), .B2(G2105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n907));
  AOI22_X1  g482(.A1(G142), .A2(new_n464), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n902), .A2(new_n908), .A3(new_n826), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n826), .B1(new_n902), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n897), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n827), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n902), .A2(new_n908), .A3(new_n826), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n639), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n895), .A2(new_n896), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n896), .B1(new_n895), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n879), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n895), .A2(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT101), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n895), .A2(new_n916), .A3(new_n896), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT102), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n895), .A2(new_n916), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G160), .B(new_n647), .ZN(new_n927));
  XNOR2_X1  g502(.A(G162), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(KEYINPUT103), .A3(new_n928), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n928), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n921), .A2(new_n922), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n931), .A2(KEYINPUT104), .A3(new_n932), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g516(.A(new_n869), .B(new_n633), .ZN(new_n942));
  NAND2_X1  g517(.A1(G299), .A2(new_n626), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n618), .A2(new_n623), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT105), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g521(.A1(G299), .A2(new_n626), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n942), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(G288), .ZN(new_n958));
  NOR3_X1   g533(.A1(G288), .A2(new_n603), .A3(new_n606), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(G303), .A2(new_n599), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n519), .B(KEYINPUT73), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n530), .B(new_n531), .ZN(new_n964));
  AOI21_X1  g539(.A(G305), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n960), .A3(KEYINPUT106), .ZN(new_n967));
  NAND2_X1  g542(.A1(G303), .A2(new_n599), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n607), .A2(new_n807), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(new_n959), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n964), .A3(G305), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n957), .B(new_n975), .ZN(new_n976));
  MUX2_X1   g551(.A(new_n866), .B(new_n976), .S(G868), .Z(G295));
  MUX2_X1   g552(.A(new_n866), .B(new_n976), .S(G868), .Z(G331));
  AOI21_X1  g553(.A(KEYINPUT77), .B1(new_n551), .B2(new_n555), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n558), .A2(new_n554), .A3(new_n557), .ZN(new_n980));
  OAI21_X1  g555(.A(G168), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n556), .A2(G286), .A3(new_n559), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n869), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n863), .A2(new_n981), .A3(new_n868), .A4(new_n982), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT108), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n869), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n953), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  INV_X1    g565(.A(new_n948), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n984), .A3(new_n985), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n989), .B2(new_n992), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n966), .A2(new_n973), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n989), .A3(new_n992), .ZN(new_n997));
  INV_X1    g572(.A(G37), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n951), .B1(new_n943), .B2(new_n944), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n948), .B2(new_n951), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n984), .A2(new_n985), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n986), .A2(new_n988), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n948), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n1008), .B2(new_n974), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n948), .B1(new_n986), .B2(new_n988), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT110), .B(new_n974), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1002), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT43), .B1(new_n996), .B2(new_n999), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n1002), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(KEYINPUT44), .B2(new_n1021), .ZN(G397));
  AOI21_X1  g597(.A(G1384), .B1(new_n889), .B2(new_n489), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(KEYINPUT45), .ZN(new_n1024));
  AND2_X1   g599(.A1(G160), .A2(G40), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1996), .ZN(new_n1027));
  INV_X1    g602(.A(new_n766), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n1029), .B(KEYINPUT111), .Z(new_n1030));
  INV_X1    g605(.A(G2067), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n723), .B(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT112), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1026), .A2(G1996), .A3(new_n766), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1026), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n826), .A2(new_n829), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n826), .A2(new_n829), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n607), .B(G1986), .Z(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1023), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1384), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n496), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT50), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1048), .A3(new_n1025), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(G1956), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n623), .B(KEYINPUT57), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1025), .B1(new_n1053), .B2(new_n1047), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1024), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1052), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(new_n709), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1025), .A2(new_n1023), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(G2067), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT118), .B1(new_n1063), .B2(new_n626), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(KEYINPUT118), .A3(new_n626), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1059), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1055), .A2(new_n1027), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1068), .A2(KEYINPUT119), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n567), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1060), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1058), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n618), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n618), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1086), .A2(new_n1087), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1067), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1062), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(G1976), .B2(new_n807), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT113), .B(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1093), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G305), .A2(G1981), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n599), .A2(new_n815), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT49), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1092), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  AOI21_X1  g682(.A(G2090), .B1(new_n1049), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1107), .B2(new_n1049), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1055), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n802), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G303), .A2(G8), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1118), .ZN(new_n1120));
  INV_X1    g695(.A(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1050), .A2(new_n703), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1106), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1055), .A2(G1966), .B1(G2084), .B2(new_n1049), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G168), .A2(new_n1121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(G8), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1127), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT51), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n1135), .C1(new_n1126), .C2(G286), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1110), .B2(G2078), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1050), .A2(G1961), .ZN(new_n1140));
  INV_X1    g715(.A(G2078), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1055), .A2(KEYINPUT53), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G171), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1139), .A2(G301), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1146), .A2(new_n1147), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  AND4_X1   g724(.A1(KEYINPUT123), .A2(new_n1144), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1125), .B(new_n1137), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1091), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1131), .A2(G286), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1106), .A2(new_n1124), .A3(new_n1119), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1106), .A2(new_n1124), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1153), .B(KEYINPUT63), .C1(new_n1120), .C2(new_n1123), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1144), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1130), .A2(new_n1162), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1125), .A4(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1100), .B(KEYINPUT116), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(G288), .A2(G1976), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1092), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1124), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n1106), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1159), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1043), .B1(new_n1152), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n720), .A2(new_n1031), .A3(new_n722), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1026), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1026), .A2(G1996), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT124), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1032), .A2(new_n1028), .ZN(new_n1181));
  OAI221_X1 g756(.A(new_n1180), .B1(KEYINPUT46), .B2(new_n1178), .C1(new_n1026), .C2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1041), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1026), .A2(G290), .A3(G1986), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT48), .Z(new_n1187));
  AOI211_X1 g762(.A(new_n1177), .B(new_n1184), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1174), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g764(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n696), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n938), .B2(new_n939), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1193), .A2(new_n1194), .A3(new_n1020), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1193), .B2(new_n1020), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1195), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1020), .ZN(G225));
endmodule


