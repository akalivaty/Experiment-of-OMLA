//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G143), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  OAI21_X1  g010(.A(G128), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT64), .A2(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(G146), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n195), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n196), .A3(G128), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT11), .A2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT11), .A2(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G137), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(G134), .A2(G137), .ZN(new_n211));
  OAI211_X1 g025(.A(G131), .B(new_n211), .C1(new_n209), .C2(G134), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n195), .B1(new_n214), .B2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n215), .A2(new_n216), .B1(new_n194), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n205), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT11), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G137), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n205), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n210), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n219), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n219), .B2(new_n229), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n213), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(G116), .B(G119), .Z(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n219), .A2(new_n229), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n213), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n204), .A2(new_n210), .A3(new_n212), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n219), .A2(new_n229), .A3(new_n230), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n245), .B2(new_n239), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n237), .B1(new_n246), .B2(new_n236), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT67), .A2(G237), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT67), .A2(G237), .ZN(new_n250));
  AOI21_X1  g064(.A(G953), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n213), .A2(new_n238), .ZN(new_n259));
  INV_X1    g073(.A(new_n236), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT28), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n236), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n245), .A2(new_n260), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n262), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n257), .B(new_n258), .C1(new_n256), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n233), .A2(new_n236), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n261), .B1(new_n271), .B2(KEYINPUT28), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n256), .A2(new_n258), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G472), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n247), .B2(new_n255), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n240), .B1(new_n233), .B2(KEYINPUT30), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n265), .B(new_n255), .C1(new_n280), .C2(new_n260), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT31), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n247), .A2(new_n284), .A3(new_n255), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n267), .A2(new_n256), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n277), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n246), .A2(new_n236), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(new_n278), .A3(new_n265), .A4(new_n255), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n284), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n286), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n277), .B(new_n289), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n276), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  MUX2_X1   g113(.A(new_n204), .B(new_n219), .S(G125), .Z(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT83), .B(G224), .ZN(new_n301));
  INV_X1    g115(.A(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(KEYINPUT7), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n234), .A2(new_n235), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n308), .A2(KEYINPUT5), .A3(G119), .ZN(new_n309));
  XNOR2_X1  g123(.A(G116), .B(G119), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(KEYINPUT5), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(G113), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT3), .A2(G107), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT3), .A2(G107), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(G104), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT74), .A2(G104), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT74), .A2(G104), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(G104), .A2(G107), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(G101), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n312), .B(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(G110), .B(G122), .Z(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT8), .Z(new_n330));
  AOI22_X1  g144(.A1(new_n304), .A2(new_n305), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n334), .A3(new_n326), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n312), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT80), .ZN(new_n337));
  INV_X1    g151(.A(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n314), .A2(G104), .ZN(new_n339));
  INV_X1    g153(.A(new_n313), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(KEYINPUT74), .A2(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT74), .A2(G104), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n314), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G101), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(G101), .C1(new_n341), .C2(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(new_n236), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n333), .A2(new_n350), .A3(new_n312), .A4(new_n335), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n337), .A2(new_n338), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n300), .A2(KEYINPUT7), .A3(new_n303), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n306), .A2(new_n331), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n337), .A2(new_n349), .A3(new_n351), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT82), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n329), .B(KEYINPUT81), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n355), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n352), .A2(new_n356), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n300), .B(new_n303), .Z(new_n363));
  OAI211_X1 g177(.A(new_n299), .B(new_n354), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G210), .B1(G237), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(new_n361), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n363), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n299), .A3(new_n365), .A4(new_n354), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(KEYINPUT85), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT79), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n364), .A2(new_n378), .A3(new_n366), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n375), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n249), .A2(new_n250), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G214), .A3(new_n302), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n199), .A2(new_n200), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n251), .A2(new_n188), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n208), .ZN(new_n388));
  OR2_X1    g202(.A1(G125), .A2(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(G125), .A2(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n190), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n384), .A2(KEYINPUT18), .A3(G131), .A4(new_n385), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n389), .B2(new_n390), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(KEYINPUT16), .A3(G140), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n389), .B(new_n390), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(new_n190), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n384), .A2(G131), .A3(new_n385), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G131), .B1(new_n384), .B2(new_n385), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n408), .B1(new_n400), .B2(new_n407), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n394), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n416), .B(G104), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT71), .B1(new_n399), .B2(G146), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT71), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n190), .C1(new_n396), .C2(new_n398), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n400), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n411), .A2(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n386), .A2(new_n208), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n410), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n424), .B(new_n425), .C1(new_n427), .C2(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n417), .A3(new_n394), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G475), .ZN(new_n431));
  AND4_X1   g245(.A1(KEYINPUT20), .A2(new_n430), .A3(new_n431), .A4(new_n299), .ZN(new_n432));
  AOI21_X1  g246(.A(G475), .B1(new_n419), .B2(new_n429), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT20), .B1(new_n433), .B2(new_n299), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n440));
  OAI21_X1  g254(.A(G478), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT9), .B(G234), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G217), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n443), .A2(new_n444), .A3(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n214), .A2(G128), .ZN(new_n446));
  INV_X1    g260(.A(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G143), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(KEYINPUT13), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n449), .B(G134), .C1(KEYINPUT13), .C2(new_n446), .ZN(new_n450));
  XNOR2_X1  g264(.A(G116), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n317), .ZN(new_n452));
  INV_X1    g266(.A(G134), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n453), .A3(new_n448), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n317), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n308), .A2(KEYINPUT14), .A3(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n451), .ZN(new_n458));
  OAI211_X1 g272(.A(G107), .B(new_n457), .C1(new_n458), .C2(KEYINPUT14), .ZN(new_n459));
  INV_X1    g273(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n453), .B1(new_n446), .B2(new_n448), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n456), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n445), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n462), .A3(new_n445), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n269), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n441), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n465), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n441), .C1(new_n469), .C2(new_n463), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n436), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n441), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n469), .A2(new_n463), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n269), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT89), .A3(new_n470), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G952), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n302), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(G234), .B2(G237), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT21), .B(G898), .Z(new_n484));
  NAND2_X1  g298(.A1(G234), .A2(G237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n269), .A2(G953), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n428), .A2(new_n394), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n417), .ZN(new_n490));
  OAI21_X1  g304(.A(G475), .B1(new_n490), .B2(G902), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n435), .A2(new_n477), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G221), .B1(new_n443), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(G469), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G140), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n302), .A2(G227), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n327), .A2(new_n204), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n201), .A2(new_n202), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n196), .B1(new_n383), .B2(new_n190), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n447), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n332), .B1(new_n501), .B2(new_n203), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n229), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n228), .A2(new_n210), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT76), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n447), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n203), .B1(new_n510), .B2(new_n215), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n327), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n332), .A2(new_n198), .A3(new_n203), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n507), .A3(new_n229), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n333), .A2(KEYINPUT10), .A3(new_n204), .A4(new_n335), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n346), .A2(new_n348), .A3(new_n219), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n505), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n497), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n346), .A2(new_n348), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n523), .A2(new_n219), .B1(new_n517), .B2(new_n512), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n505), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n497), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT77), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n514), .A2(new_n507), .A3(new_n229), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n507), .B1(new_n514), .B2(new_n229), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n497), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n521), .A2(new_n497), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n518), .A2(new_n520), .ZN(new_n536));
  INV_X1    g350(.A(new_n519), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n229), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n494), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n526), .B1(new_n515), .B2(new_n509), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n497), .B1(new_n538), .B2(new_n521), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n494), .B(new_n467), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n494), .A2(new_n299), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n493), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT78), .B(new_n493), .C1(new_n541), .C2(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n492), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n444), .B1(new_n467), .B2(G234), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n302), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(new_n222), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n557));
  INV_X1    g371(.A(G119), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(G128), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n447), .A2(KEYINPUT23), .A3(G119), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n560), .C1(G119), .C2(new_n447), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G110), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G119), .B(G128), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n423), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n391), .A2(new_n190), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n561), .A2(G110), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n400), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n568), .B2(new_n572), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n556), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n568), .A2(new_n572), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n573), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n555), .A3(new_n575), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n581), .A3(new_n467), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n582), .A2(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT73), .B1(new_n582), .B2(new_n584), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n553), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n553), .A2(G902), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n578), .A2(new_n581), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n298), .A2(new_n380), .A3(new_n552), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n550), .A2(new_n551), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n467), .B1(new_n294), .B2(new_n295), .ZN(new_n597));
  AOI22_X1  g411(.A1(G472), .A2(new_n597), .B1(new_n288), .B2(new_n289), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n595), .A2(new_n596), .A3(new_n592), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n591), .B1(new_n550), .B2(new_n551), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n595), .B1(new_n600), .B2(new_n598), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n364), .A2(new_n366), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n371), .B2(new_n372), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n365), .B1(new_n604), .B2(new_n354), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n376), .B(new_n488), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(KEYINPUT93), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(KEYINPUT93), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n474), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n474), .A2(KEYINPUT93), .A3(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(G478), .A3(new_n467), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n474), .A2(new_n269), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(G478), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n435), .A2(new_n491), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NOR3_X1   g435(.A1(new_n606), .A2(new_n477), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n602), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT94), .B(KEYINPUT35), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NAND3_X1  g440(.A1(new_n568), .A2(KEYINPUT36), .A3(new_n572), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n578), .A2(new_n581), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(KEYINPUT36), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n589), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n588), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n380), .A2(new_n552), .A3(new_n598), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G110), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(new_n376), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n367), .B2(new_n374), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n637), .A2(new_n631), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n435), .A2(new_n491), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT96), .B(G900), .Z(new_n640));
  OR2_X1    g454(.A1(new_n486), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n483), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n477), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n298), .A2(new_n638), .A3(new_n644), .A4(new_n596), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NAND2_X1  g460(.A1(new_n375), .A2(new_n379), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n631), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n477), .B1(new_n435), .B2(new_n491), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n649), .A2(new_n376), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n642), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n596), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT40), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT32), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n296), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n291), .A2(new_n293), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n271), .A2(new_n256), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n299), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT98), .ZN(new_n667));
  OR3_X1    g481(.A1(new_n652), .A2(new_n655), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n383), .ZN(G45));
  INV_X1    g483(.A(new_n642), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n617), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n298), .A2(new_n638), .A3(new_n671), .A4(new_n596), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI21_X1  g487(.A(new_n591), .B1(new_n658), .B2(new_n276), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n535), .A2(new_n516), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n538), .A2(new_n521), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n497), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n467), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(new_n493), .A3(new_n544), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n618), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n622), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  AND3_X1   g500(.A1(new_n637), .A2(new_n631), .A3(new_n680), .ZN(new_n687));
  INV_X1    g501(.A(new_n492), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n298), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  INV_X1    g504(.A(new_n680), .ZN(new_n691));
  INV_X1    g505(.A(new_n651), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n606), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n269), .B1(new_n283), .B2(new_n287), .ZN(new_n695));
  INV_X1    g509(.A(G472), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n597), .A2(KEYINPUT100), .A3(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n285), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n272), .A2(new_n255), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n294), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n289), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT99), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n701), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n283), .A2(new_n285), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT99), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n289), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n693), .A2(new_n592), .A3(new_n699), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND4_X1  g525(.A1(new_n687), .A2(new_n699), .A3(new_n709), .A4(new_n671), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  AOI21_X1  g527(.A(new_n636), .B1(new_n375), .B2(new_n379), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n298), .A2(new_n592), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n533), .A2(G469), .A3(new_n539), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n544), .A2(new_n546), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g537(.A(new_n493), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n715), .A2(new_n671), .A3(new_n718), .A4(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n298), .A2(new_n592), .A3(new_n714), .A4(new_n725), .ZN(new_n727));
  INV_X1    g541(.A(new_n671), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n716), .B(new_n717), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  NAND3_X1  g545(.A1(new_n715), .A2(new_n644), .A3(new_n725), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND3_X1  g547(.A1(new_n533), .A2(KEYINPUT45), .A3(new_n539), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT103), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n494), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n528), .A2(new_n540), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n546), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n544), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n493), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n714), .B(KEYINPUT104), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n653), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n639), .A2(new_n615), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n598), .A3(new_n650), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT44), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  NAND2_X1  g568(.A1(new_n745), .A2(KEYINPUT47), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n298), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n714), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n728), .A3(new_n592), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  AND2_X1   g576(.A1(new_n679), .A2(new_n544), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT49), .Z(new_n764));
  NAND3_X1  g578(.A1(new_n639), .A2(new_n615), .A3(new_n377), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n764), .A2(new_n591), .A3(new_n724), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n667), .A3(new_n648), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n750), .A2(new_n483), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n699), .A2(new_n709), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n592), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n648), .A2(new_n636), .A3(new_n680), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT111), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n777), .A2(KEYINPUT111), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n776), .B2(new_n778), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n763), .A2(new_n724), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n755), .A2(new_n757), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n771), .A2(new_n746), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n759), .A2(new_n691), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n592), .A2(new_n667), .A3(new_n482), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n615), .A2(new_n616), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n769), .A2(new_n787), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n631), .A3(new_n770), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n768), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n793), .B(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n783), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n755), .A2(KEYINPUT113), .A3(new_n757), .A4(new_n782), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n784), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n800), .A3(KEYINPUT51), .A4(new_n781), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n791), .A2(new_n674), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n637), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n771), .A2(new_n805), .A3(new_n691), .ZN(new_n806));
  INV_X1    g620(.A(new_n617), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n481), .B(new_n806), .C1(new_n807), .C2(new_n788), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n794), .A2(new_n801), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n699), .A2(new_n709), .A3(new_n671), .A4(new_n725), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n616), .A2(new_n471), .A3(new_n468), .A4(new_n670), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n298), .A2(new_n596), .A3(new_n812), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n650), .B(new_n759), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n727), .A2(new_n477), .A3(new_n643), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n814), .A2(KEYINPUT106), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT106), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n631), .A3(new_n714), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n819), .B2(new_n732), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n593), .A2(new_n689), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n380), .A2(new_n488), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n617), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n602), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n674), .B(new_n680), .C1(new_n622), .C2(new_n618), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n632), .A3(new_n710), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT105), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n468), .A2(new_n471), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n616), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n380), .A2(KEYINPUT105), .A3(new_n488), .A4(new_n830), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n602), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n730), .A2(new_n825), .A3(new_n827), .A4(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n651), .B(new_n376), .C1(new_n605), .C2(new_n603), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n631), .A2(new_n670), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n666), .A2(new_n837), .A3(new_n725), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n712), .A2(new_n839), .A3(new_n645), .A4(new_n672), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n821), .A2(new_n835), .A3(KEYINPUT53), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT108), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n825), .A2(new_n827), .A3(new_n834), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n730), .A3(new_n842), .ZN(new_n848));
  INV_X1    g662(.A(new_n820), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n819), .A2(new_n817), .A3(new_n732), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n846), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n825), .A2(new_n730), .A3(new_n827), .A4(new_n834), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n712), .A2(new_n645), .A3(new_n672), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n841), .A3(new_n839), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT108), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n844), .A2(new_n845), .A3(new_n852), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n855), .A2(KEYINPUT107), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n846), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n858), .A2(new_n863), .A3(new_n821), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n858), .B2(new_n821), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n810), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n866), .A3(new_n810), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n809), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(G952), .A2(G953), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n767), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT115), .B(new_n767), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(G75));
  NAND3_X1  g690(.A1(new_n844), .A2(new_n852), .A3(new_n860), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n269), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n366), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n371), .B(new_n363), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n879), .B2(new_n880), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n302), .A2(G952), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G51));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n877), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n877), .B2(KEYINPUT54), .ZN(new_n889));
  INV_X1    g703(.A(new_n861), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n545), .B(KEYINPUT57), .Z(new_n892));
  OAI21_X1  g706(.A(new_n677), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n739), .B(KEYINPUT117), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n885), .B1(new_n893), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n430), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n885), .ZN(G60));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n902));
  INV_X1    g716(.A(new_n885), .ZN(new_n903));
  INV_X1    g717(.A(new_n612), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n861), .A2(new_n810), .A3(new_n866), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n867), .ZN(new_n911));
  INV_X1    g725(.A(new_n906), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n612), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n902), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n889), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n877), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n861), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n885), .B1(new_n917), .B2(new_n907), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n868), .A2(new_n869), .A3(new_n912), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(KEYINPUT118), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(G63));
  XNOR2_X1  g736(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n444), .A2(new_n299), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n877), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n885), .B1(new_n926), .B2(new_n628), .ZN(new_n927));
  INV_X1    g741(.A(new_n629), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n926), .ZN(new_n929));
  XOR2_X1   g743(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G66));
  AOI21_X1  g745(.A(new_n302), .B1(new_n484), .B2(new_n301), .ZN(new_n932));
  INV_X1    g746(.A(new_n847), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n302), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n362), .B1(G898), .B2(new_n302), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(G69));
  AOI21_X1  g750(.A(new_n654), .B1(new_n617), .B2(new_n831), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n715), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n748), .B2(new_n752), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n761), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n854), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n668), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(new_n947));
  OAI21_X1  g761(.A(new_n302), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n280), .B(KEYINPUT121), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n403), .A2(new_n406), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(G900), .A2(G953), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n753), .A2(new_n854), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n745), .A2(new_n674), .A3(new_n653), .A4(new_n837), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n758), .B2(new_n760), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n958), .A2(KEYINPUT125), .B1(new_n726), .B2(new_n729), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n957), .A2(new_n960), .A3(new_n732), .A4(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n955), .B(new_n956), .C1(new_n962), .C2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n948), .A2(KEYINPUT124), .A3(new_n951), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n954), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n302), .B1(G227), .B2(G900), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n864), .B2(new_n865), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n257), .B(KEYINPUT126), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n659), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT127), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n969), .B1(new_n962), .B2(new_n933), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n247), .A3(new_n256), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n942), .A2(new_n947), .A3(new_n933), .ZN(new_n976));
  INV_X1    g790(.A(new_n969), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n248), .B(new_n255), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AND4_X1   g792(.A1(new_n903), .A2(new_n973), .A3(new_n975), .A4(new_n978), .ZN(G57));
endmodule


