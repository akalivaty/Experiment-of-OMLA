//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n191), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n188), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n193), .A2(G143), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n197), .A2(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n190), .B2(new_n207), .ZN(new_n208));
  AND4_X1   g022(.A1(new_n206), .A2(new_n207), .A3(new_n194), .A4(new_n196), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n202), .B(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G224), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n211), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G110), .B(G122), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT2), .B(G113), .Z(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT68), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G107), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n230), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT81), .A2(G107), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n232), .B(new_n234), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  AOI21_X1  g055(.A(G101), .B1(new_n233), .B2(G107), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n232), .B(new_n242), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n245), .A3(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n229), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n218), .ZN(new_n248));
  OAI21_X1  g062(.A(G113), .B1(new_n221), .B2(KEYINPUT5), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(KEYINPUT5), .B2(new_n217), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT81), .A2(G107), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT81), .A2(G107), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n254), .A2(new_n255), .B1(KEYINPUT3), .B2(new_n231), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n233), .B1(new_n252), .B2(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n231), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n256), .A2(new_n242), .B1(new_n258), .B2(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  AOI211_X1 g074(.A(KEYINPUT6), .B(new_n215), .C1(new_n247), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n244), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n227), .A3(new_n228), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n215), .B(new_n260), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n247), .A2(KEYINPUT88), .A3(new_n215), .A4(new_n260), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n215), .B1(new_n247), .B2(new_n260), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n214), .B(new_n261), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n266), .A2(new_n267), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n211), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n249), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(new_n224), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n249), .A2(new_n277), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n218), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n259), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n215), .B(KEYINPUT8), .Z(new_n284));
  AOI21_X1  g098(.A(G104), .B1(new_n236), .B2(new_n237), .ZN(new_n285));
  INV_X1    g099(.A(new_n231), .ZN(new_n286));
  OAI21_X1  g100(.A(G101), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n243), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n284), .B1(new_n251), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n276), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n201), .A2(new_n210), .A3(KEYINPUT90), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n190), .B2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n207), .A2(new_n194), .A3(new_n196), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n190), .A2(new_n206), .A3(new_n207), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT90), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n202), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n275), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n291), .A2(new_n299), .A3(KEYINPUT91), .A4(new_n275), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n273), .B1(new_n274), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n272), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n268), .A2(new_n271), .ZN(new_n309));
  INV_X1    g123(.A(new_n261), .ZN(new_n310));
  INV_X1    g124(.A(new_n214), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n290), .A2(new_n302), .A3(new_n303), .ZN(new_n313));
  AOI21_X1  g127(.A(G902), .B1(new_n313), .B2(new_n268), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n306), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n187), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT14), .ZN(new_n317));
  INV_X1    g131(.A(G122), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n317), .A2(new_n318), .A3(G116), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G122), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n230), .B(new_n319), .C1(new_n317), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n254), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n195), .A2(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n203), .A2(G143), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n322), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT13), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT13), .B1(new_n195), .B2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n323), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(KEYINPUT98), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n337), .A3(new_n323), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n325), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n222), .A2(G122), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n318), .A2(G116), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n340), .A2(new_n341), .B1(new_n253), .B2(new_n252), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n326), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT99), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n332), .B1(new_n203), .B2(G143), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n203), .A2(G143), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT98), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n333), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n338), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G134), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n327), .B1(new_n342), .B2(new_n322), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT99), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n331), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n331), .B(new_n360), .C1(new_n346), .C2(new_n354), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n273), .ZN(new_n363));
  INV_X1    g177(.A(G478), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT15), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(new_n365), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n212), .A3(G214), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G143), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n195), .A2(KEYINPUT92), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G237), .A2(G953), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n375), .A2(G214), .B1(new_n371), .B2(G143), .ZN(new_n376));
  OAI21_X1  g190(.A(G131), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n372), .ZN(new_n378));
  INV_X1    g192(.A(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT92), .B(G143), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n378), .B(new_n379), .C1(new_n370), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n202), .A2(G140), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(KEYINPUT16), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT76), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G146), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT19), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT19), .B1(new_n384), .B2(new_n385), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n193), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n382), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT18), .B(G131), .C1(new_n374), .C2(new_n376), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n384), .A2(new_n385), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n384), .A2(new_n385), .A3(new_n193), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n374), .A2(new_n376), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT93), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n379), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n378), .B(new_n407), .C1(new_n370), .C2(new_n380), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n381), .A2(new_n409), .A3(KEYINPUT93), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n404), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n398), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n377), .A2(new_n413), .A3(new_n381), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT94), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n193), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n418));
  OR3_X1    g232(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT76), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n193), .B1(new_n420), .B2(new_n387), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n377), .A2(new_n381), .A3(new_n423), .A4(new_n413), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n377), .A2(new_n413), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n415), .A2(new_n422), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n408), .A2(new_n410), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n399), .A3(new_n403), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n397), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n412), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n397), .B1(new_n426), .B2(new_n428), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n434), .A2(KEYINPUT95), .A3(new_n412), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(KEYINPUT20), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n431), .A2(KEYINPUT95), .A3(new_n437), .A4(new_n432), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(KEYINPUT100), .A2(G952), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT100), .A2(G952), .ZN(new_n442));
  AOI21_X1  g256(.A(G953), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G234), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n369), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n273), .B(new_n212), .C1(G234), .C2(G237), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(G898), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n397), .A2(KEYINPUT97), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n429), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n429), .A2(new_n451), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n273), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT96), .B(G475), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n368), .A2(new_n439), .A3(new_n450), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n316), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n297), .B2(new_n288), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n259), .A2(KEYINPUT10), .A3(new_n462), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT69), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT69), .B1(new_n192), .B2(new_n199), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n244), .B(new_n246), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G137), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G134), .ZN(new_n471));
  NOR2_X1   g285(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n325), .A2(G137), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n325), .A2(G137), .ZN(new_n477));
  AND2_X1   g291(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n478), .B2(new_n472), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n471), .A2(new_n474), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n379), .A3(new_n476), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n465), .A2(new_n466), .A3(new_n469), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n259), .B2(new_n462), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n297), .A2(new_n288), .A3(KEYINPUT85), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n461), .A3(new_n463), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT12), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT84), .B1(new_n480), .B2(new_n483), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n493), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n489), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(G110), .B(G140), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT80), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n212), .A2(G227), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n489), .A2(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n484), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G469), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT86), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n500), .A2(new_n505), .B1(new_n509), .B2(new_n507), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(G469), .C1(new_n515), .C2(G902), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n498), .A2(new_n499), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n489), .A2(new_n504), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT87), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n507), .B(new_n520), .C1(new_n498), .C2(new_n499), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n509), .A2(new_n489), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n505), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n512), .A3(new_n273), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n516), .A3(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n458), .A2(new_n459), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT77), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G137), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT78), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n220), .B2(G128), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n535), .B(new_n536), .C1(G119), .C2(new_n203), .ZN(new_n537));
  XNOR2_X1  g351(.A(G119), .B(G128), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT24), .B(G110), .Z(new_n539));
  AOI22_X1  g353(.A1(new_n537), .A2(G110), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n417), .B2(new_n421), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n537), .A2(G110), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n391), .A2(new_n542), .A3(new_n402), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n544), .A2(new_n531), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n273), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n546), .A4(new_n273), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n357), .B1(G234), .B2(new_n273), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n551), .B(KEYINPUT75), .Z(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(G902), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n546), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT79), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n484), .B1(new_n467), .B2(new_n468), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n471), .A2(new_n476), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G131), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n483), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n462), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(KEYINPUT30), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT70), .A4(KEYINPUT30), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n200), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n462), .A2(new_n563), .B1(new_n484), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT67), .B1(new_n571), .B2(KEYINPUT30), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT67), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n483), .A2(new_n562), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n297), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n200), .B1(new_n483), .B2(new_n480), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n573), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n579), .A3(new_n229), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n227), .A2(new_n228), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n560), .A2(new_n581), .A3(new_n564), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n375), .A2(G210), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT27), .Z(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT26), .B(G101), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT31), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n580), .A2(KEYINPUT31), .A3(new_n588), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT72), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT28), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n229), .B1(new_n576), .B2(new_n577), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n582), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT69), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n190), .A2(new_n189), .A3(new_n191), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n188), .B1(new_n197), .B2(new_n198), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT69), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(new_n483), .B2(new_n480), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n603), .B2(new_n576), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n560), .A2(KEYINPUT71), .A3(new_n564), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n581), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n596), .B1(new_n594), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n587), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n593), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n560), .A2(new_n564), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n229), .B1(new_n610), .B2(new_n597), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT28), .B1(new_n611), .B2(new_n605), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT72), .B(new_n587), .C1(new_n612), .C2(new_n596), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n591), .A2(new_n592), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT32), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n606), .A2(new_n594), .ZN(new_n618));
  INV_X1    g432(.A(new_n596), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT72), .B1(new_n620), .B2(new_n587), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n607), .A2(new_n593), .A3(new_n608), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n580), .A2(KEYINPUT31), .A3(new_n588), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT31), .B1(new_n580), .B2(new_n588), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT32), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n615), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n617), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n567), .A2(new_n568), .B1(new_n572), .B2(new_n578), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n583), .B1(new_n629), .B2(new_n229), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT73), .B1(new_n630), .B2(new_n608), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n580), .A2(new_n582), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT73), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n587), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT29), .B1(new_n607), .B2(new_n608), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n581), .B1(new_n560), .B2(new_n564), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT28), .B1(new_n583), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n608), .A2(KEYINPUT29), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n618), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT74), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n640), .A2(new_n641), .A3(new_n273), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n640), .B2(new_n273), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n559), .B1(new_n628), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n527), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G101), .ZN(G3));
  OAI21_X1  g463(.A(G472), .B1(new_n614), .B2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n625), .A2(new_n615), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n559), .ZN(new_n653));
  INV_X1    g467(.A(new_n459), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n489), .B(new_n504), .C1(new_n498), .C2(new_n499), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(KEYINPUT87), .B1(new_n505), .B2(new_n522), .ZN(new_n656));
  AOI21_X1  g470(.A(G902), .B1(new_n656), .B2(new_n521), .ZN(new_n657));
  OAI21_X1  g471(.A(G469), .B1(new_n515), .B2(G902), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n512), .A2(new_n657), .B1(new_n658), .B2(KEYINPUT86), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n654), .B1(new_n659), .B2(new_n516), .ZN(new_n660));
  INV_X1    g474(.A(new_n187), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n307), .B1(new_n272), .B2(new_n305), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n312), .A2(new_n314), .A3(new_n306), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n450), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n429), .A2(new_n430), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  INV_X1    g481(.A(new_n412), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n669), .A2(new_n437), .B1(new_n431), .B2(new_n432), .ZN(new_n670));
  AND4_X1   g484(.A1(KEYINPUT95), .A2(new_n431), .A3(new_n437), .A4(new_n432), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n456), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n363), .A2(new_n364), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n345), .B1(new_n339), .B2(new_n344), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n352), .A2(KEYINPUT99), .A3(new_n353), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n330), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n360), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n330), .B(new_n358), .C1(new_n674), .C2(new_n675), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n678), .A3(KEYINPUT33), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n361), .A2(KEYINPUT102), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n358), .A2(KEYINPUT102), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n355), .A2(KEYINPUT101), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n681), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n679), .B1(KEYINPUT33), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n273), .A2(G478), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n673), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n672), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n665), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n653), .A2(new_n660), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT34), .B(G104), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G6));
  AOI21_X1  g508(.A(new_n437), .B1(new_n431), .B2(new_n432), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n431), .A2(new_n437), .A3(new_n432), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n368), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n456), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n665), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n653), .A2(new_n660), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT35), .B(G107), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G9));
  NOR2_X1   g519(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n544), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n554), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n553), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n652), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n527), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT37), .B(G110), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G12));
  NAND2_X1  g528(.A1(new_n628), .A2(new_n646), .ZN(new_n715));
  INV_X1    g529(.A(new_n445), .ZN(new_n716));
  INV_X1    g530(.A(G900), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n717), .B2(new_n446), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n700), .A2(new_n699), .A3(new_n456), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n664), .A2(new_n709), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n715), .A2(new_n660), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT105), .B(G128), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G30));
  NAND2_X1  g539(.A1(new_n526), .A2(new_n459), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n718), .B(KEYINPUT39), .Z(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OR3_X1    g542(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT40), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT108), .B1(new_n726), .B2(new_n728), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n587), .B1(new_n580), .B2(new_n582), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n583), .A2(new_n637), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n273), .B1(new_n736), .B2(new_n608), .ZN(new_n737));
  OAI21_X1  g551(.A(G472), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT106), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n628), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n662), .A2(new_n663), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT38), .ZN(new_n742));
  INV_X1    g556(.A(new_n672), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n743), .A2(new_n661), .A3(new_n709), .A4(new_n368), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n740), .A2(KEYINPUT107), .A3(new_n742), .A4(new_n744), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n733), .A2(new_n734), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n195), .ZN(G45));
  NAND3_X1  g565(.A1(new_n672), .A2(new_n689), .A3(new_n719), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n672), .A2(new_n689), .A3(new_n754), .A4(new_n719), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n715), .A3(new_n660), .A4(new_n722), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G146), .ZN(G48));
  NAND2_X1  g572(.A1(new_n524), .A2(new_n273), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(G469), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n459), .A3(new_n525), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n647), .A2(new_n691), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT41), .B(G113), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT110), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n763), .B(new_n765), .ZN(G15));
  NAND3_X1  g580(.A1(new_n647), .A2(new_n702), .A3(new_n762), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G116), .ZN(G18));
  NAND4_X1  g582(.A1(new_n760), .A2(new_n459), .A3(new_n664), .A4(new_n525), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n457), .A2(new_n710), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n715), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G119), .ZN(G21));
  INV_X1    g587(.A(new_n559), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n618), .A2(new_n638), .ZN(new_n775));
  OAI22_X1  g589(.A1(new_n623), .A2(new_n624), .B1(new_n608), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n615), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n591), .A2(new_n592), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n609), .A2(new_n613), .ZN(new_n779));
  AOI21_X1  g593(.A(G902), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(G472), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n774), .B(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n650), .A2(KEYINPUT111), .A3(new_n774), .A4(new_n777), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n368), .B1(new_n456), .B2(new_n439), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n664), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n761), .A2(new_n788), .A3(new_n449), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G122), .ZN(G24));
  NAND2_X1  g605(.A1(new_n753), .A2(new_n755), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n709), .B(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n792), .A2(new_n769), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n202), .ZN(G27));
  INV_X1    g609(.A(new_n489), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n493), .A2(new_n497), .ZN(new_n797));
  INV_X1    g611(.A(new_n496), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n510), .B1(new_n801), .B2(new_n504), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n512), .B1(new_n802), .B2(new_n273), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n657), .B2(new_n512), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n662), .A2(new_n663), .A3(new_n459), .A4(new_n187), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n756), .A2(new_n715), .A3(new_n774), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n647), .A2(new_n756), .A3(KEYINPUT42), .A4(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G131), .ZN(G33));
  NAND3_X1  g626(.A1(new_n647), .A2(new_n720), .A3(new_n806), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  NAND2_X1  g628(.A1(new_n515), .A2(KEYINPUT45), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(G469), .B1(new_n515), .B2(KEYINPUT45), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(G469), .A2(G902), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n820), .A2(new_n821), .B1(new_n512), .B2(new_n657), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(KEYINPUT46), .A3(new_n819), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n654), .B(new_n728), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n662), .A2(new_n663), .A3(new_n187), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT112), .Z(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n743), .A2(new_n828), .A3(new_n689), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n743), .B2(new_n689), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n710), .B1(new_n650), .B2(new_n651), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n827), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n652), .A2(new_n709), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT44), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n824), .B(new_n826), .C1(new_n834), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G137), .ZN(G39));
  AOI21_X1  g654(.A(new_n654), .B1(new_n822), .B2(new_n823), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n617), .A2(new_n627), .B1(new_n645), .B2(G472), .ZN(new_n844));
  INV_X1    g658(.A(new_n825), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n756), .A2(new_n844), .A3(new_n559), .A4(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT113), .B(G140), .Z(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(G42));
  AND2_X1   g663(.A1(new_n760), .A2(new_n525), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT114), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n743), .A2(new_n689), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n774), .A2(new_n459), .A3(new_n187), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n740), .A2(new_n742), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n718), .A2(new_n654), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n708), .A2(new_n553), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT115), .B1(new_n804), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n788), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n525), .A2(new_n658), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  INV_X1    g679(.A(new_n861), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n740), .A2(new_n862), .A3(new_n863), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n793), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n756), .A2(new_n770), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n757), .A2(new_n723), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n859), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n647), .B(new_n762), .C1(new_n691), .C2(new_n702), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n368), .A2(new_n439), .A3(new_n456), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n743), .B2(new_n689), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n665), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n653), .A2(new_n881), .A3(new_n660), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n878), .A2(new_n772), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n527), .B1(new_n647), .B2(new_n711), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(new_n790), .ZN(new_n885));
  INV_X1    g699(.A(new_n699), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n709), .A2(new_n368), .A3(new_n456), .A4(new_n719), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n825), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n715), .A2(new_n660), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n756), .A2(new_n869), .A3(new_n806), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n813), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n883), .A2(new_n885), .A3(new_n811), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n844), .A2(new_n726), .A3(new_n721), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n788), .B1(new_n628), .B2(new_n739), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT115), .B(new_n861), .C1(new_n525), .C2(new_n658), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n897), .A2(new_n756), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n794), .B1(new_n897), .B2(new_n720), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT52), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n874), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n896), .B1(new_n906), .B2(new_n892), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n894), .A2(new_n895), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n878), .A2(new_n772), .A3(new_n882), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n884), .A2(new_n790), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n813), .A2(new_n889), .A3(new_n890), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n809), .B2(new_n810), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n905), .A2(KEYINPUT53), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT117), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n893), .A2(new_n916), .A3(KEYINPUT53), .A4(new_n905), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n892), .B1(new_n875), .B2(new_n876), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n915), .B(new_n917), .C1(KEYINPUT53), .C2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n908), .B1(KEYINPUT54), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n850), .A2(new_n845), .A3(new_n459), .A4(new_n716), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(new_n836), .ZN(new_n922));
  INV_X1    g736(.A(new_n647), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT48), .Z(new_n925));
  AND3_X1   g739(.A1(new_n786), .A2(new_n716), .A3(new_n832), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n770), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT118), .ZN(new_n928));
  INV_X1    g742(.A(new_n443), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n921), .A2(new_n559), .A3(new_n740), .ZN(new_n930));
  INV_X1    g744(.A(new_n690), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n851), .A2(new_n654), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n843), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n826), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n742), .A2(new_n761), .A3(new_n187), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n926), .A2(KEYINPUT50), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT50), .B1(new_n926), .B2(new_n939), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT51), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n922), .A2(new_n793), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n672), .A2(new_n689), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n930), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n938), .A2(new_n942), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n940), .B2(new_n941), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n936), .B1(new_n843), .B2(new_n934), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT51), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n933), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT119), .B1(new_n920), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n915), .A2(new_n917), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n918), .A2(KEYINPUT53), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT54), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n894), .A2(new_n895), .A3(new_n907), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(KEYINPUT119), .A3(new_n956), .A4(new_n951), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT120), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n858), .B1(new_n952), .B2(new_n960), .ZN(G75));
  NOR2_X1   g775(.A1(new_n212), .A2(G952), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n273), .B1(new_n894), .B2(new_n907), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT56), .B1(new_n964), .B2(G210), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n261), .B1(new_n268), .B2(new_n271), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n311), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(new_n272), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT55), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n965), .B2(new_n970), .ZN(G51));
  XNOR2_X1  g786(.A(new_n818), .B(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n819), .B(KEYINPUT57), .Z(new_n977));
  AOI21_X1  g791(.A(new_n895), .B1(new_n894), .B2(new_n907), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n908), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n524), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n962), .B1(new_n976), .B2(new_n980), .ZN(G54));
  INV_X1    g795(.A(new_n431), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT58), .ZN(new_n983));
  INV_X1    g797(.A(G475), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n896), .B(new_n892), .C1(new_n875), .C2(new_n876), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT53), .B1(new_n893), .B2(new_n905), .ZN(new_n989));
  OAI211_X1 g803(.A(G902), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT123), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n964), .A2(new_n992), .A3(new_n987), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n273), .B(new_n986), .C1(new_n894), .C2(new_n907), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n963), .B1(new_n995), .B2(new_n431), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT124), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n964), .A2(new_n985), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n962), .B1(new_n998), .B2(new_n982), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT124), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(new_n1000), .A3(new_n991), .A4(new_n993), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1001), .ZN(G60));
  INV_X1    g816(.A(new_n687), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n955), .A2(new_n956), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G478), .A2(G902), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT59), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1003), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1003), .B(new_n1006), .C1(new_n908), .C2(new_n978), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n963), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1007), .A2(new_n1009), .ZN(G63));
  NAND2_X1  g824(.A1(G217), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT60), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n894), .B2(new_n907), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n545), .A2(new_n546), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1013), .A2(new_n707), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n963), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT61), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1016), .A2(KEYINPUT61), .A3(new_n963), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(G66));
  INV_X1    g836(.A(G224), .ZN(new_n1023));
  OAI21_X1  g837(.A(G953), .B1(new_n447), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n911), .B2(G953), .ZN(new_n1025));
  INV_X1    g839(.A(G898), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n966), .B1(new_n1026), .B2(G953), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT125), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1025), .B(new_n1028), .ZN(G69));
  AOI21_X1  g843(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n392), .A2(new_n393), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n629), .B(new_n1031), .Z(new_n1032));
  NOR2_X1   g846(.A1(new_n880), .A2(new_n825), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n729), .A2(new_n647), .A3(new_n731), .A4(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n839), .A2(KEYINPUT126), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n826), .B1(new_n838), .B2(new_n834), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n841), .A2(new_n727), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n903), .A2(new_n757), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT62), .B1(new_n750), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT62), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1042), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n749), .A2(new_n734), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n733), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n1041), .A2(new_n1043), .A3(new_n847), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1032), .B1(new_n1048), .B2(new_n212), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT127), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(G900), .A2(G953), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n824), .A2(new_n647), .A3(new_n863), .ZN(new_n1054));
  AND3_X1   g868(.A1(new_n1054), .A2(new_n811), .A3(new_n813), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n847), .A2(new_n839), .A3(new_n1045), .A4(new_n1055), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n1032), .B(new_n1053), .C1(new_n1056), .C2(G953), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1057), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1030), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1048), .A2(new_n212), .ZN(new_n1060));
  OAI21_X1  g874(.A(KEYINPUT127), .B1(new_n1060), .B2(new_n1032), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1030), .ZN(new_n1062));
  NAND4_X1  g876(.A1(new_n1061), .A2(new_n1062), .A3(new_n1051), .A4(new_n1057), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1059), .A2(new_n1063), .ZN(G72));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  NAND3_X1  g880(.A1(new_n631), .A2(new_n589), .A3(new_n634), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n919), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(new_n911), .ZN(new_n1069));
  OAI21_X1  g883(.A(new_n1066), .B1(new_n1056), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n632), .A2(new_n608), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n1068), .A2(new_n1072), .A3(new_n963), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1066), .B1(new_n1048), .B2(new_n1069), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1073), .B1(new_n735), .B2(new_n1074), .ZN(G57));
endmodule


