//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n467), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n463), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT67), .Z(new_n487));
  AOI211_X1 g062(.A(new_n483), .B(new_n487), .C1(G136), .C2(new_n469), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n468), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  AOI211_X1 g066(.A(G2105), .B(new_n489), .C1(KEYINPUT68), .C2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n492), .A2(new_n472), .A3(new_n467), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n485), .B2(G126), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT69), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n506), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  XNOR2_X1  g088(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n503), .B2(new_n504), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n507), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT5), .B(G543), .Z(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n505), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n518), .A2(new_n528), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n507), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n519), .A2(new_n524), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G52), .A3(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(G90), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n527), .A2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n507), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n530), .A2(G81), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G860), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g123(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n549));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(new_n530), .ZN(new_n553));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n553), .A2(new_n554), .B1(new_n507), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n526), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n519), .A2(new_n524), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT74), .A4(new_n560), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n561), .B2(new_n562), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n572));
  NOR2_X1   g147(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n558), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g150(.A(KEYINPUT77), .B(new_n573), .C1(new_n567), .C2(new_n570), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n557), .B1(new_n575), .B2(new_n576), .ZN(G299));
  NOR2_X1   g152(.A1(G171), .A2(KEYINPUT78), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(G301));
  OR2_X1    g157(.A1(new_n501), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(G651), .A2(new_n583), .B1(new_n530), .B2(G87), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n527), .A2(KEYINPUT79), .A3(G49), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT79), .B1(new_n527), .B2(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n589), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n529), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n501), .A2(KEYINPUT81), .A3(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n501), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n505), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n527), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n507), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n530), .A2(G85), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n530), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT10), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n527), .A2(G54), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(G66), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(G66), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n501), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G79), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n526), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G651), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n609), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n618), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g194(.A(new_n618), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT75), .B1(new_n569), .B2(new_n564), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n574), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT77), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n573), .B1(new_n567), .B2(new_n570), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n558), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n556), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n621), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(new_n618), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n545), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n618), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n638));
  XNOR2_X1  g213(.A(G323), .B(new_n638), .ZN(G282));
  NAND2_X1  g214(.A1(new_n469), .A2(G135), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT84), .Z(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n642), .A2(KEYINPUT85), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(KEYINPUT85), .B2(new_n642), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n484), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n657));
  XOR2_X1   g232(.A(KEYINPUT15), .B(G2435), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XOR2_X1   g234(.A(G2427), .B(G2430), .Z(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n698), .B(new_n699), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(new_n703), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n685), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n704), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n703), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(new_n684), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n469), .A2(G131), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT88), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(G107), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G2105), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n485), .B2(G119), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n715), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G16), .A2(G24), .ZN(new_n726));
  INV_X1    g301(.A(G290), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT89), .B(G1986), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G22), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G166), .B2(new_n731), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1971), .ZN(new_n734));
  MUX2_X1   g309(.A(G6), .B(G305), .S(G16), .Z(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT32), .B(G1981), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G23), .B(new_n587), .S(G16), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT33), .B(G1976), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n737), .B(new_n740), .C1(new_n735), .C2(new_n736), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n725), .B(new_n730), .C1(new_n741), .C2(KEYINPUT34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(KEYINPUT34), .B2(new_n741), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT36), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n731), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT23), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n628), .B2(new_n731), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n731), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n731), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT97), .Z(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  INV_X1    g329(.A(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT24), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n479), .B2(new_n714), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n469), .A2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n485), .A2(G129), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n767), .A2(new_n768), .B1(new_n477), .B2(G105), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G129), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(new_n484), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G141), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n468), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT92), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  MUX2_X1   g353(.A(KEYINPUT93), .B(new_n761), .S(new_n778), .Z(new_n779));
  OAI21_X1  g354(.A(new_n759), .B1(new_n760), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n714), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n714), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT29), .Z(new_n784));
  INV_X1    g359(.A(G2090), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G4), .A2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT90), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n618), .B2(new_n731), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n649), .A2(new_n714), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT95), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n752), .A2(new_n753), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n731), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n731), .B2(G21), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT94), .B(G1966), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT96), .Z(new_n800));
  NAND4_X1  g375(.A1(new_n786), .A2(new_n794), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n797), .A2(new_n798), .B1(new_n754), .B2(new_n758), .ZN(new_n802));
  INV_X1    g377(.A(G28), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT30), .ZN(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n803), .B2(KEYINPUT30), .ZN(new_n805));
  OR2_X1    g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  NAND2_X1  g381(.A1(KEYINPUT31), .A2(G11), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G19), .B(new_n545), .S(G16), .Z(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G1341), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n714), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  INV_X1    g388(.A(G140), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n468), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT91), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G116), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n485), .B2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n813), .B1(new_n822), .B2(new_n714), .ZN(new_n823));
  INV_X1    g398(.A(G2067), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n714), .A2(G27), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G164), .B2(new_n714), .ZN(new_n827));
  INV_X1    g402(.A(G2078), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n714), .A2(G33), .ZN(new_n830));
  NAND2_X1  g405(.A1(G115), .A2(G2104), .ZN(new_n831));
  INV_X1    g406(.A(G127), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n473), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n834));
  NAND2_X1  g409(.A1(G103), .A2(G2104), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(G2105), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n833), .A2(G2105), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n469), .A2(G139), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n830), .B1(new_n841), .B2(new_n714), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G2072), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G1341), .B2(new_n809), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n811), .A2(new_n825), .A3(new_n829), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n779), .A2(new_n760), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n784), .B2(new_n785), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n801), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n744), .A2(new_n749), .A3(new_n781), .A4(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  NAND2_X1  g425(.A1(new_n631), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n529), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n855), .A2(G651), .B1(new_n530), .B2(G93), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n527), .A2(G55), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n545), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n852), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n546), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(new_n649), .B(new_n479), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(G162), .Z(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n722), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n776), .A2(G164), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n495), .A2(new_n499), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n770), .A3(new_n775), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n822), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n841), .B2(KEYINPUT100), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n841), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n821), .A3(new_n874), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n878), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n876), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n871), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n469), .A2(G142), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n485), .A2(G130), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n466), .A2(G118), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(new_n653), .Z(new_n890));
  INV_X1    g465(.A(new_n880), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n821), .B1(new_n872), .B2(new_n874), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n878), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n722), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n884), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n890), .B1(new_n884), .B2(new_n895), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n870), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(new_n897), .A3(new_n869), .A4(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g481(.A1(new_n858), .A2(new_n634), .ZN(new_n907));
  NAND2_X1  g482(.A1(G299), .A2(new_n618), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n631), .B(new_n557), .C1(new_n575), .C2(new_n576), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n628), .A2(new_n631), .ZN(new_n912));
  AOI211_X1 g487(.A(new_n556), .B(new_n618), .C1(new_n625), .C2(new_n627), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n915), .A3(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n859), .B(KEYINPUT103), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n636), .ZN(new_n919));
  MUX2_X1   g494(.A(new_n911), .B(new_n917), .S(new_n919), .Z(new_n920));
  XNOR2_X1  g495(.A(G166), .B(G305), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n587), .B(new_n727), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n926), .B(new_n927), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n920), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n907), .B1(new_n929), .B2(new_n634), .ZN(G295));
  OAI21_X1  g505(.A(new_n907), .B1(new_n929), .B2(new_n634), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n908), .A2(new_n909), .A3(new_n934), .A4(new_n915), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n914), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G168), .B1(new_n578), .B2(new_n581), .ZN(new_n937));
  NAND2_X1  g512(.A1(G286), .A2(new_n579), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n937), .A2(new_n859), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n859), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n932), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n910), .A2(new_n941), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n936), .A2(new_n932), .A3(new_n941), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n926), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n908), .A2(new_n915), .A3(new_n909), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n915), .B1(new_n908), .B2(new_n909), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n941), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n943), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n926), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n904), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n939), .A2(new_n940), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n914), .B2(new_n916), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT106), .B1(new_n958), .B2(new_n943), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n950), .A2(new_n960), .A3(new_n951), .ZN(new_n961));
  INV_X1    g536(.A(new_n926), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n954), .B(KEYINPUT44), .C1(new_n956), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n952), .A2(new_n955), .A3(new_n904), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n945), .A2(new_n942), .A3(new_n943), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n926), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n964), .A3(new_n952), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n970), .C2(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n966), .B1(new_n975), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  XNOR2_X1  g553(.A(G305), .B(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(KEYINPUT49), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(KEYINPUT49), .ZN(new_n981));
  NAND2_X1  g556(.A1(G160), .A2(G40), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n873), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n588), .A2(new_n989), .A3(new_n590), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n587), .A2(new_n989), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n990), .A2(new_n987), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n992), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT52), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT113), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n982), .B1(new_n1001), .B2(new_n984), .ZN(new_n1002));
  INV_X1    g577(.A(new_n984), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1006));
  AND2_X1   g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1005), .A2(G1971), .B1(G2090), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1000), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n999), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n997), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n984), .A2(new_n1001), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n1016), .B2(new_n982), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1002), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(G2078), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1017), .A2(new_n1019), .A3(new_n1004), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1009), .A2(new_n753), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1002), .A2(new_n828), .A3(new_n1004), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1020), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(KEYINPUT121), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(KEYINPUT121), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(new_n1023), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G301), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1014), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1017), .A2(new_n1004), .A3(new_n1019), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n798), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n754), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1036), .B2(G286), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1038));
  AOI21_X1  g613(.A(G168), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1031), .A2(new_n1038), .A3(KEYINPUT62), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1011), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1013), .B1(new_n1010), .B2(G8), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n996), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G286), .A2(new_n986), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1036), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1044), .B(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT63), .B1(new_n1051), .B2(new_n1014), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n980), .A2(new_n981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n989), .A3(new_n591), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(G1981), .B2(G305), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n987), .A2(new_n1055), .B1(new_n997), .B2(new_n1042), .ZN(new_n1056));
  AND4_X1   g631(.A1(new_n1041), .A2(new_n1050), .A3(new_n1052), .A4(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1014), .A2(new_n1030), .A3(KEYINPUT62), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1009), .A2(new_n790), .B1(new_n985), .B2(new_n824), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n631), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n631), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1059), .A2(new_n631), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1002), .A2(new_n1066), .A3(new_n1004), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n982), .B2(new_n984), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n545), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1002), .A2(new_n1004), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1034), .B2(G1956), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n628), .A2(KEYINPUT57), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n626), .B2(new_n556), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1076), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(G299), .B2(new_n1078), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1005), .A2(new_n1074), .B1(new_n1009), .B2(new_n748), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(KEYINPUT61), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1082), .A2(new_n1085), .A3(KEYINPUT120), .A4(KEYINPUT61), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1073), .A2(new_n1088), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1083), .A2(new_n1084), .B1(new_n618), .B2(new_n1059), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1094), .A2(new_n1085), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT54), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1023), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1009), .A2(KEYINPUT122), .A3(new_n753), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(G2078), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1005), .A2(KEYINPUT53), .A3(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n579), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1044), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1101), .A2(new_n1107), .A3(G301), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT54), .B1(new_n1110), .B2(new_n1030), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1058), .B1(new_n1099), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1057), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1015), .A2(new_n982), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(G1996), .A3(new_n776), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1066), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n776), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT111), .Z(new_n1121));
  XNOR2_X1  g696(.A(new_n821), .B(G2067), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1118), .B(new_n1121), .C1(new_n1116), .C2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n722), .A2(new_n724), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n722), .A2(new_n724), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G290), .A2(G1986), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(KEYINPUT110), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G290), .A2(G1986), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1129), .B(new_n1130), .Z(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1116), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT46), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT124), .Z(new_n1136));
  OAI21_X1  g711(.A(new_n777), .B1(new_n1134), .B2(G1996), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1116), .B1(new_n1122), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT47), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT126), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1143));
  XNOR2_X1  g718(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1140), .B1(new_n1127), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(G2067), .B2(new_n821), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1116), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1133), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g724(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1151));
  AOI21_X1  g725(.A(new_n1151), .B1(new_n708), .B2(new_n711), .ZN(new_n1152));
  NAND2_X1  g726(.A1(new_n905), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g727(.A(new_n1153), .ZN(new_n1154));
  AND3_X1   g728(.A1(new_n973), .A2(KEYINPUT127), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g729(.A(KEYINPUT127), .B1(new_n973), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1156), .ZN(G308));
  NAND2_X1  g731(.A1(new_n973), .A2(new_n1154), .ZN(new_n1158));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n973), .A2(new_n1154), .A3(KEYINPUT127), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1161), .ZN(G225));
endmodule


