

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(n663), .ZN(n681) );
  OR2_X1 U554 ( .A1(KEYINPUT33), .A2(n712), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n738), .A2(n745), .ZN(n739) );
  OR2_X1 U556 ( .A1(n634), .A2(n973), .ZN(n633) );
  XNOR2_X1 U557 ( .A(n671), .B(KEYINPUT99), .ZN(n673) );
  NAND2_X1 U558 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U559 ( .A(n689), .B(n688), .ZN(n697) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  AND2_X1 U561 ( .A1(n716), .A2(n521), .ZN(n520) );
  OR2_X1 U562 ( .A1(n715), .A2(n714), .ZN(n521) );
  NOR2_X1 U563 ( .A1(n714), .A2(n710), .ZN(n522) );
  OR2_X1 U564 ( .A1(n706), .A2(n705), .ZN(n523) );
  INV_X1 U565 ( .A(G8), .ZN(n668) );
  OR2_X1 U566 ( .A1(n690), .A2(n668), .ZN(n669) );
  OR2_X1 U567 ( .A1(n693), .A2(n669), .ZN(n670) );
  XNOR2_X1 U568 ( .A(n633), .B(KEYINPUT98), .ZN(n655) );
  INV_X1 U569 ( .A(G168), .ZN(n672) );
  AND2_X1 U570 ( .A1(n673), .A2(n672), .ZN(n676) );
  XNOR2_X1 U571 ( .A(n662), .B(KEYINPUT29), .ZN(n667) );
  INV_X1 U572 ( .A(KEYINPUT32), .ZN(n688) );
  NAND2_X1 U573 ( .A1(n697), .A2(n696), .ZN(n708) );
  NAND2_X1 U574 ( .A1(G8), .A2(n681), .ZN(n714) );
  INV_X1 U575 ( .A(G40), .ZN(n588) );
  AND2_X2 U576 ( .A1(n527), .A2(G2104), .ZN(n885) );
  NOR2_X1 U577 ( .A1(G651), .A2(n568), .ZN(n800) );
  XOR2_X1 U578 ( .A(KEYINPUT17), .B(n524), .Z(n582) );
  BUF_X1 U579 ( .A(n582), .Z(n884) );
  NAND2_X1 U580 ( .A1(G138), .A2(n884), .ZN(n526) );
  INV_X1 U581 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U582 ( .A1(G102), .A2(n885), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n532) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U585 ( .A1(n888), .A2(G114), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n527), .A2(G2104), .ZN(n528) );
  XNOR2_X1 U587 ( .A(n528), .B(KEYINPUT64), .ZN(n584) );
  BUF_X1 U588 ( .A(n584), .Z(n889) );
  NAND2_X1 U589 ( .A1(G126), .A2(n889), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n532), .A2(n531), .ZN(G164) );
  INV_X1 U592 ( .A(G651), .ZN(n536) );
  NOR2_X1 U593 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n533), .Z(n796) );
  NAND2_X1 U595 ( .A1(G64), .A2(n796), .ZN(n535) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n568) );
  NAND2_X1 U597 ( .A1(G52), .A2(n800), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n797) );
  NAND2_X1 U600 ( .A1(G90), .A2(n797), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n568), .A2(n536), .ZN(n801) );
  NAND2_X1 U602 ( .A1(G77), .A2(n801), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(G171) );
  NAND2_X1 U606 ( .A1(n797), .A2(G89), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G76), .A2(n801), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n796), .A2(G63), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT72), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G51), .A2(n800), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G88), .A2(n797), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G75), .A2(n801), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G62), .A2(n796), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT79), .B(n555), .Z(n557) );
  NAND2_X1 U624 ( .A1(n800), .A2(G50), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(G166) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  NAND2_X1 U628 ( .A1(G61), .A2(n796), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G86), .A2(n797), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n801), .A2(G73), .ZN(n562) );
  XOR2_X1 U632 ( .A(KEYINPUT2), .B(n562), .Z(n563) );
  NOR2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT78), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G48), .A2(n800), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(G305) );
  NAND2_X1 U637 ( .A1(G49), .A2(n800), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G87), .A2(n568), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U640 ( .A1(n796), .A2(n571), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n572) );
  XOR2_X1 U642 ( .A(KEYINPUT77), .B(n572), .Z(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U644 ( .A1(G60), .A2(n796), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G47), .A2(n800), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(n577), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G85), .A2(n797), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G72), .A2(n801), .ZN(n578) );
  AND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(G290) );
  NAND2_X1 U652 ( .A1(G137), .A2(n582), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT66), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n584), .A2(G125), .ZN(n585) );
  XOR2_X1 U655 ( .A(n585), .B(KEYINPUT65), .Z(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n779) );
  NOR2_X1 U657 ( .A1(n779), .A2(n588), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n888), .A2(G113), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G101), .A2(n885), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT23), .B(n589), .Z(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n780) );
  INV_X1 U662 ( .A(n780), .ZN(n592) );
  AND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT84), .ZN(n619) );
  INV_X1 U665 ( .A(n619), .ZN(n595) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n620) );
  NOR2_X1 U667 ( .A1(n595), .A2(n620), .ZN(n752) );
  XNOR2_X1 U668 ( .A(KEYINPUT37), .B(G2067), .ZN(n750) );
  XNOR2_X1 U669 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n888), .A2(G116), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G128), .A2(n889), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT35), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n600), .B(n599), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n885), .A2(G104), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT85), .B(n601), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n884), .A2(G140), .ZN(n602) );
  XOR2_X1 U678 ( .A(KEYINPUT86), .B(n602), .Z(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U680 ( .A(KEYINPUT34), .B(n605), .Z(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U682 ( .A(KEYINPUT36), .B(n608), .ZN(n904) );
  OR2_X1 U683 ( .A1(n750), .A2(n904), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT89), .ZN(n928) );
  NAND2_X1 U685 ( .A1(n752), .A2(n928), .ZN(n748) );
  NAND2_X1 U686 ( .A1(G56), .A2(n796), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(n610), .Z(n616) );
  NAND2_X1 U688 ( .A1(n797), .A2(G81), .ZN(n611) );
  XNOR2_X1 U689 ( .A(n611), .B(KEYINPUT12), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G68), .A2(n801), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U692 ( .A(KEYINPUT13), .B(n614), .Z(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n800), .A2(G43), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n988) );
  AND2_X2 U696 ( .A1(n620), .A2(n619), .ZN(n663) );
  NAND2_X1 U697 ( .A1(G1996), .A2(n663), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT26), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G1341), .A2(n681), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U701 ( .A(KEYINPUT96), .B(n624), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n988), .A2(n625), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G66), .A2(n796), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G92), .A2(n797), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G54), .A2(n800), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G79), .A2(n801), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U710 ( .A(KEYINPUT15), .B(n632), .Z(n973) );
  NAND2_X1 U711 ( .A1(n634), .A2(n973), .ZN(n639) );
  INV_X1 U712 ( .A(G2067), .ZN(n950) );
  NOR2_X1 U713 ( .A1(n681), .A2(n950), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n635), .B(KEYINPUT97), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n681), .A2(G1348), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n653) );
  NAND2_X1 U718 ( .A1(G91), .A2(n797), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G78), .A2(n801), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(KEYINPUT68), .B(n642), .ZN(n646) );
  NAND2_X1 U722 ( .A1(G65), .A2(n796), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G53), .A2(n800), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT69), .B(n647), .Z(n972) );
  XOR2_X1 U727 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n649) );
  NAND2_X1 U728 ( .A1(G2072), .A2(n663), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U730 ( .A(G1956), .ZN(n1000) );
  NOR2_X1 U731 ( .A1(n663), .A2(n1000), .ZN(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n657) );
  NOR2_X1 U733 ( .A1(n972), .A2(n657), .ZN(n652) );
  XOR2_X1 U734 ( .A(n652), .B(KEYINPUT28), .Z(n656) );
  AND2_X1 U735 ( .A1(n653), .A2(n656), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n661) );
  INV_X1 U737 ( .A(n656), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n972), .A2(n657), .ZN(n658) );
  OR2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NOR2_X1 U741 ( .A1(n681), .A2(n956), .ZN(n665) );
  INV_X1 U742 ( .A(G1961), .ZN(n1009) );
  NOR2_X1 U743 ( .A1(n663), .A2(n1009), .ZN(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n674) );
  NAND2_X1 U745 ( .A1(G171), .A2(n674), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n680) );
  NOR2_X1 U747 ( .A1(G1966), .A2(n714), .ZN(n693) );
  NOR2_X1 U748 ( .A1(G2084), .A2(n681), .ZN(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT30), .B(n670), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G171), .A2(n674), .ZN(n675) );
  NOR2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n678) );
  INV_X1 U752 ( .A(KEYINPUT31), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U754 ( .A1(n680), .A2(n679), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n691), .A2(G286), .ZN(n687) );
  NOR2_X1 U756 ( .A1(G1971), .A2(n714), .ZN(n683) );
  NOR2_X1 U757 ( .A1(G2090), .A2(n681), .ZN(n682) );
  NOR2_X1 U758 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n684), .A2(G303), .ZN(n685) );
  OR2_X1 U760 ( .A1(n668), .A2(n685), .ZN(n686) );
  NAND2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U762 ( .A1(G8), .A2(n690), .ZN(n695) );
  INV_X1 U763 ( .A(n691), .ZN(n692) );
  NOR2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U767 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n708), .A2(n699), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n700), .A2(n714), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT101), .ZN(n706) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XOR2_X1 U772 ( .A(n702), .B(KEYINPUT24), .Z(n703) );
  NOR2_X1 U773 ( .A1(n714), .A2(n703), .ZN(n704) );
  XNOR2_X1 U774 ( .A(n704), .B(KEYINPUT94), .ZN(n705) );
  NAND2_X1 U775 ( .A1(n748), .A2(n523), .ZN(n718) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n713) );
  NOR2_X1 U777 ( .A1(G1971), .A2(G303), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n713), .A2(n707), .ZN(n978) );
  NAND2_X1 U779 ( .A1(n708), .A2(n978), .ZN(n709) );
  XNOR2_X1 U780 ( .A(n709), .B(KEYINPUT100), .ZN(n711) );
  NAND2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U782 ( .A(n977), .ZN(n710) );
  AND2_X1 U783 ( .A1(n711), .A2(n522), .ZN(n712) );
  XOR2_X1 U784 ( .A(G1981), .B(G305), .Z(n969) );
  AND2_X1 U785 ( .A1(n969), .A2(n748), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n713), .A2(KEYINPUT33), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n519), .A2(n520), .ZN(n717) );
  AND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n738) );
  NAND2_X1 U789 ( .A1(G95), .A2(n885), .ZN(n719) );
  XNOR2_X1 U790 ( .A(n719), .B(KEYINPUT90), .ZN(n726) );
  NAND2_X1 U791 ( .A1(n888), .A2(G107), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G119), .A2(n889), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U794 ( .A1(G131), .A2(n884), .ZN(n722) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n722), .ZN(n723) );
  NOR2_X1 U796 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n898) );
  NAND2_X1 U798 ( .A1(G1991), .A2(n898), .ZN(n736) );
  XOR2_X1 U799 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n728) );
  NAND2_X1 U800 ( .A1(G105), .A2(n885), .ZN(n727) );
  XNOR2_X1 U801 ( .A(n728), .B(n727), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G141), .A2(n884), .ZN(n730) );
  NAND2_X1 U803 ( .A1(G117), .A2(n888), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U806 ( .A1(G129), .A2(n889), .ZN(n733) );
  NAND2_X1 U807 ( .A1(n734), .A2(n733), .ZN(n897) );
  NAND2_X1 U808 ( .A1(G1996), .A2(n897), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n921) );
  NAND2_X1 U810 ( .A1(n921), .A2(n752), .ZN(n737) );
  XNOR2_X1 U811 ( .A(n737), .B(KEYINPUT93), .ZN(n745) );
  XNOR2_X1 U812 ( .A(n739), .B(KEYINPUT102), .ZN(n741) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U814 ( .A1(n984), .A2(n752), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n755) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n897), .ZN(n742) );
  XOR2_X1 U817 ( .A(KEYINPUT103), .B(n742), .Z(n918) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n898), .ZN(n924) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n924), .A2(n743), .ZN(n744) );
  NOR2_X1 U821 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U822 ( .A1(n918), .A2(n746), .ZN(n747) );
  XNOR2_X1 U823 ( .A(n747), .B(KEYINPUT39), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n904), .A2(n750), .ZN(n932) );
  NAND2_X1 U826 ( .A1(n751), .A2(n932), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U830 ( .A(G2443), .B(G2435), .ZN(n766) );
  XOR2_X1 U831 ( .A(G2427), .B(KEYINPUT105), .Z(n758) );
  XNOR2_X1 U832 ( .A(G2454), .B(G2430), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n758), .B(n757), .ZN(n762) );
  XOR2_X1 U834 ( .A(KEYINPUT104), .B(G2446), .Z(n760) );
  XNOR2_X1 U835 ( .A(G1348), .B(G1341), .ZN(n759) );
  XNOR2_X1 U836 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U837 ( .A(n762), .B(n761), .Z(n764) );
  XNOR2_X1 U838 ( .A(G2451), .B(G2438), .ZN(n763) );
  XNOR2_X1 U839 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U840 ( .A(n766), .B(n765), .ZN(n767) );
  AND2_X1 U841 ( .A1(n767), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U843 ( .A1(G111), .A2(n888), .ZN(n776) );
  NAND2_X1 U844 ( .A1(G135), .A2(n884), .ZN(n769) );
  NAND2_X1 U845 ( .A1(G99), .A2(n885), .ZN(n768) );
  NAND2_X1 U846 ( .A1(n769), .A2(n768), .ZN(n774) );
  XOR2_X1 U847 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n771) );
  NAND2_X1 U848 ( .A1(G123), .A2(n889), .ZN(n770) );
  XNOR2_X1 U849 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U850 ( .A(KEYINPUT74), .B(n772), .Z(n773) );
  NOR2_X1 U851 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U852 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n777), .B(KEYINPUT76), .ZN(n922) );
  XNOR2_X1 U854 ( .A(n922), .B(G2096), .ZN(n778) );
  OR2_X1 U855 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G57), .ZN(G237) );
  NOR2_X1 U859 ( .A1(n779), .A2(n780), .ZN(G160) );
  XOR2_X1 U860 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n782) );
  NAND2_X1 U861 ( .A1(G7), .A2(G661), .ZN(n781) );
  XNOR2_X1 U862 ( .A(n782), .B(n781), .ZN(G223) );
  INV_X1 U863 ( .A(G223), .ZN(n836) );
  NAND2_X1 U864 ( .A1(n836), .A2(G567), .ZN(n783) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n783), .Z(G234) );
  INV_X1 U866 ( .A(G860), .ZN(n788) );
  OR2_X1 U867 ( .A1(n988), .A2(n788), .ZN(G153) );
  INV_X1 U868 ( .A(G171), .ZN(G301) );
  NAND2_X1 U869 ( .A1(G868), .A2(G301), .ZN(n785) );
  OR2_X1 U870 ( .A1(n973), .A2(G868), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(G284) );
  XOR2_X1 U872 ( .A(n972), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n787) );
  INV_X1 U874 ( .A(G868), .ZN(n817) );
  NOR2_X1 U875 ( .A1(G286), .A2(n817), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(G297) );
  NAND2_X1 U877 ( .A1(n788), .A2(G559), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n789), .A2(n973), .ZN(n790) );
  XNOR2_X1 U879 ( .A(n790), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U880 ( .A1(G868), .A2(n988), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G868), .A2(n973), .ZN(n791) );
  NOR2_X1 U882 ( .A1(G559), .A2(n791), .ZN(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U884 ( .A(KEYINPUT73), .B(n794), .Z(G282) );
  NAND2_X1 U885 ( .A1(n973), .A2(G559), .ZN(n813) );
  XNOR2_X1 U886 ( .A(n988), .B(n813), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n795), .A2(G860), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G93), .A2(n797), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G55), .A2(n800), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n816) );
  XOR2_X1 U895 ( .A(n806), .B(n816), .Z(G145) );
  XNOR2_X1 U896 ( .A(KEYINPUT19), .B(G290), .ZN(n807) );
  XNOR2_X1 U897 ( .A(n807), .B(G288), .ZN(n808) );
  XNOR2_X1 U898 ( .A(G299), .B(n808), .ZN(n811) );
  XNOR2_X1 U899 ( .A(n816), .B(G166), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n809), .B(n988), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n812), .B(G305), .ZN(n907) );
  XNOR2_X1 U903 ( .A(n907), .B(n813), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(G868), .ZN(n815) );
  XNOR2_X1 U905 ( .A(n815), .B(KEYINPUT80), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XOR2_X1 U911 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n822) );
  XNOR2_X1 U912 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U915 ( .A1(G69), .A2(G120), .ZN(n825) );
  NOR2_X1 U916 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U917 ( .A1(G108), .A2(n826), .ZN(n841) );
  NAND2_X1 U918 ( .A1(G567), .A2(n841), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT83), .ZN(n833) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n828) );
  XNOR2_X1 U921 ( .A(KEYINPUT22), .B(n828), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(G96), .ZN(n830) );
  NOR2_X1 U923 ( .A1(n830), .A2(G218), .ZN(n831) );
  XOR2_X1 U924 ( .A(n831), .B(KEYINPUT82), .Z(n840) );
  AND2_X1 U925 ( .A1(n840), .A2(G2106), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G319) );
  INV_X1 U927 ( .A(G319), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G483), .A2(G661), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2474), .B(G1956), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1966), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n844), .B(KEYINPUT108), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U948 ( .A(G1961), .B(G1971), .Z(n848) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1976), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U952 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U954 ( .A(G2678), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(KEYINPUT42), .B(G2090), .Z(n856) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(G2096), .B(G2100), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U963 ( .A(G2078), .B(G2084), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G227) );
  NAND2_X1 U965 ( .A1(G124), .A2(n889), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G136), .A2(n884), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT110), .B(n866), .Z(n868) );
  NAND2_X1 U970 ( .A1(n888), .A2(G112), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G100), .A2(n885), .ZN(n869) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n869), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n873) );
  XNOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n883) );
  NAND2_X1 U978 ( .A1(n888), .A2(G118), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G130), .A2(n889), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G142), .A2(n884), .ZN(n877) );
  NAND2_X1 U982 ( .A1(G106), .A2(n885), .ZN(n876) );
  NAND2_X1 U983 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  XNOR2_X1 U985 ( .A(KEYINPUT112), .B(n879), .ZN(n880) );
  NOR2_X1 U986 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U987 ( .A(n883), .B(n882), .Z(n896) );
  NAND2_X1 U988 ( .A1(G139), .A2(n884), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G103), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U991 ( .A1(n888), .A2(G115), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G127), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n935) );
  XNOR2_X1 U996 ( .A(G164), .B(n935), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n922), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G160), .B(G162), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1005 ( .A(n907), .B(G286), .Z(n909) );
  XNOR2_X1 U1006 ( .A(G171), .B(n973), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n911), .B(KEYINPUT49), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT115), .B(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT51), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1025 ( .A(KEYINPUT116), .B(n926), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT117), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT118), .B(n934), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G2072), .B(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G164), .B(G2078), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT119), .B(n938), .Z(n939) );
  XNOR2_X1 U1035 ( .A(KEYINPUT50), .B(n939), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n945), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(G1996), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(n946), .B(G32), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G1991), .B(G25), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n949), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT120), .B(n950), .Z(n951) );
  XNOR2_X1 U1048 ( .A(G26), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1051 ( .A(G27), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT53), .B(n959), .Z(n962) );
  XOR2_X1 U1054 ( .A(KEYINPUT54), .B(G34), .Z(n960) );
  XNOR2_X1 U1055 ( .A(G2084), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n966), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT122), .B(n967), .Z(n968) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n968), .ZN(n1024) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT57), .ZN(n992) );
  XNOR2_X1 U1067 ( .A(n972), .B(G1956), .ZN(n986) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n973), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT123), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G171), .B(n1009), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n982) );
  AND2_X1 U1072 ( .A1(G303), .A2(G1971), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT124), .B(n987), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1341), .B(n988), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1022) );
  INV_X1 U1083 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1084 ( .A(G1976), .B(G23), .Z(n996) );
  XOR2_X1 U1085 ( .A(G1971), .B(G22), .Z(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G24), .B(G1986), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(n999), .Z(n1016) );
  XNOR2_X1 U1090 ( .A(G20), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .Z(n1005) );
  XNOR2_X1 U1096 ( .A(G4), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1009), .B(G5), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT126), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT61), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

