

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741;

  INV_X1 U362 ( .A(KEYINPUT126), .ZN(n343) );
  NAND2_X1 U363 ( .A1(n380), .A2(n571), .ZN(n379) );
  AND2_X1 U364 ( .A1(n505), .A2(n715), .ZN(n380) );
  XNOR2_X1 U365 ( .A(n452), .B(n451), .ZN(n517) );
  XNOR2_X1 U366 ( .A(n511), .B(KEYINPUT1), .ZN(n555) );
  XNOR2_X1 U367 ( .A(n398), .B(n429), .ZN(n600) );
  NAND2_X1 U368 ( .A1(n407), .A2(n405), .ZN(n514) );
  XNOR2_X1 U369 ( .A(n463), .B(n462), .ZN(n562) );
  XNOR2_X1 U370 ( .A(n483), .B(n444), .ZN(n456) );
  INV_X1 U371 ( .A(G128), .ZN(n443) );
  XNOR2_X1 U372 ( .A(G119), .B(KEYINPUT3), .ZN(n734) );
  XNOR2_X1 U373 ( .A(KEYINPUT67), .B(G101), .ZN(n494) );
  XNOR2_X1 U374 ( .A(n372), .B(n374), .ZN(n392) );
  XNOR2_X2 U375 ( .A(n410), .B(KEYINPUT81), .ZN(n509) );
  XNOR2_X1 U376 ( .A(n344), .B(n343), .ZN(G66) );
  NAND2_X1 U377 ( .A1(n651), .A2(n687), .ZN(n344) );
  NAND2_X2 U378 ( .A1(n360), .A2(n377), .ZN(n376) );
  OR2_X2 U379 ( .A1(n693), .A2(G902), .ZN(n502) );
  INV_X1 U380 ( .A(G953), .ZN(n725) );
  BUF_X1 U381 ( .A(G128), .Z(n708) );
  XNOR2_X2 U382 ( .A(n672), .B(G146), .ZN(n496) );
  NOR2_X1 U383 ( .A1(n660), .A2(n656), .ZN(n402) );
  XNOR2_X1 U384 ( .A(n574), .B(n403), .ZN(n656) );
  XNOR2_X1 U385 ( .A(n509), .B(KEYINPUT19), .ZN(n548) );
  XNOR2_X1 U386 ( .A(G146), .B(G125), .ZN(n485) );
  XNOR2_X1 U387 ( .A(n566), .B(n565), .ZN(n660) );
  XNOR2_X2 U388 ( .A(n594), .B(KEYINPUT45), .ZN(n722) );
  XNOR2_X2 U389 ( .A(n456), .B(n412), .ZN(n672) );
  XNOR2_X1 U390 ( .A(G140), .B(G137), .ZN(n668) );
  XNOR2_X1 U391 ( .A(n364), .B(G107), .ZN(n479) );
  XNOR2_X1 U392 ( .A(G122), .B(G116), .ZN(n364) );
  AND2_X1 U393 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U394 ( .A(n570), .B(n354), .ZN(n366) );
  NAND2_X1 U395 ( .A1(n662), .A2(n489), .ZN(n452) );
  XOR2_X1 U396 ( .A(G113), .B(G116), .Z(n447) );
  NOR2_X1 U397 ( .A1(n740), .A2(n657), .ZN(n535) );
  INV_X1 U398 ( .A(KEYINPUT68), .ZN(n417) );
  XNOR2_X1 U399 ( .A(n379), .B(KEYINPUT101), .ZN(n540) );
  INV_X1 U400 ( .A(KEYINPUT8), .ZN(n413) );
  INV_X1 U401 ( .A(G110), .ZN(n421) );
  XNOR2_X1 U402 ( .A(n481), .B(n373), .ZN(n372) );
  XNOR2_X1 U403 ( .A(n397), .B(KEYINPUT39), .ZN(n547) );
  OR2_X1 U404 ( .A1(n534), .A2(n533), .ZN(n397) );
  AND2_X1 U405 ( .A1(n612), .A2(n530), .ZN(n531) );
  OR2_X1 U406 ( .A1(n648), .A2(G902), .ZN(n398) );
  INV_X1 U407 ( .A(n575), .ZN(n596) );
  INV_X1 U408 ( .A(n571), .ZN(n365) );
  AND2_X2 U409 ( .A1(n371), .A2(n381), .ZN(n692) );
  NAND2_X1 U410 ( .A1(n369), .A2(n367), .ZN(n371) );
  OR2_X1 U411 ( .A1(n387), .A2(n368), .ZN(n367) );
  NAND2_X1 U412 ( .A1(n639), .A2(n386), .ZN(n385) );
  INV_X1 U413 ( .A(KEYINPUT79), .ZN(n386) );
  XNOR2_X1 U414 ( .A(n482), .B(KEYINPUT4), .ZN(n373) );
  XNOR2_X1 U415 ( .A(n517), .B(KEYINPUT6), .ZN(n571) );
  XNOR2_X1 U416 ( .A(n496), .B(n390), .ZN(n662) );
  XNOR2_X1 U417 ( .A(n449), .B(n445), .ZN(n390) );
  AND2_X1 U418 ( .A1(n357), .A2(n349), .ZN(n673) );
  INV_X1 U419 ( .A(KEYINPUT48), .ZN(n358) );
  XOR2_X1 U420 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n453) );
  NAND2_X1 U421 ( .A1(n388), .A2(KEYINPUT2), .ZN(n387) );
  NAND2_X1 U422 ( .A1(n487), .A2(KEYINPUT79), .ZN(n388) );
  INV_X1 U423 ( .A(n385), .ZN(n368) );
  NAND2_X1 U424 ( .A1(n487), .A2(n595), .ZN(n384) );
  NAND2_X1 U425 ( .A1(n370), .A2(n722), .ZN(n369) );
  AND2_X1 U426 ( .A1(n673), .A2(n385), .ZN(n370) );
  BUF_X1 U427 ( .A(n389), .Z(n382) );
  INV_X1 U428 ( .A(KEYINPUT34), .ZN(n559) );
  XNOR2_X1 U429 ( .A(n480), .B(n479), .ZN(n393) );
  XNOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n476) );
  XNOR2_X1 U431 ( .A(n399), .B(n420), .ZN(n648) );
  XNOR2_X1 U432 ( .A(n424), .B(n419), .ZN(n399) );
  XNOR2_X1 U433 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U434 ( .A(n396), .B(n395), .ZN(n657) );
  INV_X1 U435 ( .A(KEYINPUT40), .ZN(n395) );
  INV_X1 U436 ( .A(n572), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n361), .B(n378), .ZN(n360) );
  INV_X1 U438 ( .A(KEYINPUT36), .ZN(n378) );
  INV_X1 U439 ( .A(KEYINPUT32), .ZN(n403) );
  AND2_X1 U440 ( .A1(n366), .A2(n350), .ZN(n576) );
  NAND2_X1 U441 ( .A1(n345), .A2(n362), .ZN(n715) );
  INV_X1 U442 ( .A(KEYINPUT56), .ZN(n355) );
  AND2_X1 U443 ( .A1(n363), .A2(n348), .ZN(n345) );
  AND2_X1 U444 ( .A1(n562), .A2(n503), .ZN(n346) );
  XNOR2_X1 U445 ( .A(n554), .B(KEYINPUT85), .ZN(n347) );
  OR2_X1 U446 ( .A1(n503), .A2(KEYINPUT100), .ZN(n348) );
  AND2_X1 U447 ( .A1(n741), .A2(n654), .ZN(n349) );
  AND2_X1 U448 ( .A1(n575), .A2(n517), .ZN(n350) );
  AND2_X1 U449 ( .A1(n579), .A2(n517), .ZN(n351) );
  AND2_X1 U450 ( .A1(n568), .A2(n567), .ZN(n352) );
  AND2_X1 U451 ( .A1(n503), .A2(KEYINPUT100), .ZN(n353) );
  XOR2_X1 U452 ( .A(n569), .B(KEYINPUT65), .Z(n354) );
  XNOR2_X1 U453 ( .A(n501), .B(n500), .ZN(n693) );
  INV_X1 U454 ( .A(KEYINPUT2), .ZN(n595) );
  NAND2_X1 U455 ( .A1(n684), .A2(n489), .ZN(n475) );
  XNOR2_X1 U456 ( .A(n472), .B(n473), .ZN(n684) );
  NAND2_X1 U457 ( .A1(n692), .A2(G210), .ZN(n645) );
  NAND2_X1 U458 ( .A1(n540), .A2(n509), .ZN(n361) );
  XNOR2_X1 U459 ( .A(n359), .B(n358), .ZN(n357) );
  XNOR2_X1 U460 ( .A(n376), .B(KEYINPUT80), .ZN(n375) );
  XNOR2_X1 U461 ( .A(n356), .B(n355), .ZN(G51) );
  NAND2_X1 U462 ( .A1(n647), .A2(n687), .ZN(n356) );
  NAND2_X1 U463 ( .A1(n537), .A2(n536), .ZN(n359) );
  NAND2_X1 U464 ( .A1(n353), .A2(n562), .ZN(n362) );
  OR2_X1 U465 ( .A1(n562), .A2(KEYINPUT100), .ZN(n363) );
  AND2_X1 U466 ( .A1(n366), .A2(n365), .ZN(n588) );
  NAND2_X1 U467 ( .A1(n722), .A2(n673), .ZN(n389) );
  XNOR2_X1 U468 ( .A(n486), .B(n483), .ZN(n374) );
  NAND2_X1 U469 ( .A1(n383), .A2(n384), .ZN(n381) );
  INV_X1 U470 ( .A(n376), .ZN(n658) );
  NAND2_X1 U471 ( .A1(n524), .A2(n375), .ZN(n525) );
  INV_X1 U472 ( .A(n389), .ZN(n383) );
  XNOR2_X1 U473 ( .A(n382), .B(n595), .ZN(n640) );
  NAND2_X1 U474 ( .A1(n391), .A2(n352), .ZN(n570) );
  NAND2_X1 U475 ( .A1(n607), .A2(n391), .ZN(n584) );
  XNOR2_X1 U476 ( .A(n391), .B(KEYINPUT86), .ZN(n394) );
  XNOR2_X2 U477 ( .A(n400), .B(KEYINPUT0), .ZN(n391) );
  NAND2_X1 U478 ( .A1(n641), .A2(n492), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n392), .B(n393), .ZN(n641) );
  XNOR2_X1 U480 ( .A(n393), .B(n735), .ZN(n737) );
  NAND2_X1 U481 ( .A1(n620), .A2(n394), .ZN(n560) );
  AND2_X1 U482 ( .A1(n394), .A2(n351), .ZN(n580) );
  NAND2_X1 U483 ( .A1(n547), .A2(n346), .ZN(n396) );
  NOR2_X2 U484 ( .A1(n548), .A2(n347), .ZN(n400) );
  XNOR2_X1 U485 ( .A(n401), .B(n578), .ZN(n593) );
  NAND2_X1 U486 ( .A1(n655), .A2(n402), .ZN(n401) );
  XNOR2_X2 U487 ( .A(n404), .B(KEYINPUT98), .ZN(n655) );
  NAND2_X1 U488 ( .A1(n577), .A2(n586), .ZN(n404) );
  OR2_X1 U489 ( .A1(n641), .A2(n406), .ZN(n405) );
  OR2_X1 U490 ( .A1(n492), .A2(n487), .ZN(n406) );
  NAND2_X1 U491 ( .A1(n492), .A2(n487), .ZN(n408) );
  NAND2_X1 U492 ( .A1(n514), .A2(n611), .ZN(n410) );
  AND2_X1 U493 ( .A1(n457), .A2(G217), .ZN(n411) );
  XOR2_X1 U494 ( .A(KEYINPUT4), .B(G131), .Z(n412) );
  XNOR2_X1 U495 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n608) );
  XNOR2_X1 U496 ( .A(n609), .B(n608), .ZN(n610) );
  INV_X1 U497 ( .A(KEYINPUT119), .ZN(n624) );
  INV_X1 U498 ( .A(G134), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n494), .B(G104), .ZN(n495) );
  XNOR2_X1 U500 ( .A(n624), .B(KEYINPUT52), .ZN(n625) );
  XNOR2_X1 U501 ( .A(n481), .B(n448), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n626), .B(n625), .ZN(n627) );
  INV_X1 U503 ( .A(G478), .ZN(n461) );
  XNOR2_X1 U504 ( .A(n458), .B(n411), .ZN(n459) );
  XNOR2_X1 U505 ( .A(n461), .B(KEYINPUT97), .ZN(n462) );
  INV_X1 U506 ( .A(KEYINPUT121), .ZN(n636) );
  NOR2_X1 U507 ( .A1(n562), .A2(n503), .ZN(n719) );
  XNOR2_X1 U508 ( .A(n638), .B(n637), .ZN(G75) );
  NAND2_X1 U509 ( .A1(n725), .A2(G234), .ZN(n414) );
  XNOR2_X1 U510 ( .A(n414), .B(n413), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n457), .A2(G221), .ZN(n416) );
  XNOR2_X1 U512 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n415) );
  XNOR2_X1 U513 ( .A(n416), .B(n415), .ZN(n420) );
  XNOR2_X1 U514 ( .A(n417), .B(KEYINPUT10), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n418), .B(n485), .ZN(n670) );
  INV_X1 U516 ( .A(n670), .ZN(n419) );
  XNOR2_X1 U517 ( .A(n668), .B(n421), .ZN(n499) );
  XNOR2_X1 U518 ( .A(n708), .B(G119), .ZN(n422) );
  XNOR2_X1 U519 ( .A(n422), .B(KEYINPUT87), .ZN(n423) );
  XNOR2_X1 U520 ( .A(n499), .B(n423), .ZN(n424) );
  INV_X1 U521 ( .A(KEYINPUT15), .ZN(n425) );
  XNOR2_X1 U522 ( .A(n425), .B(G902), .ZN(n487) );
  INV_X1 U523 ( .A(n487), .ZN(n639) );
  NAND2_X1 U524 ( .A1(n639), .A2(G234), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n426), .B(KEYINPUT20), .ZN(n435) );
  AND2_X1 U526 ( .A1(n435), .A2(G217), .ZN(n428) );
  XNOR2_X1 U527 ( .A(KEYINPUT76), .B(KEYINPUT25), .ZN(n427) );
  XNOR2_X1 U528 ( .A(n428), .B(n427), .ZN(n429) );
  NAND2_X1 U529 ( .A1(G234), .A2(G237), .ZN(n430) );
  XNOR2_X1 U530 ( .A(n430), .B(KEYINPUT14), .ZN(n432) );
  NAND2_X1 U531 ( .A1(G952), .A2(n432), .ZN(n628) );
  NOR2_X1 U532 ( .A1(G953), .A2(n628), .ZN(n431) );
  XNOR2_X1 U533 ( .A(n431), .B(KEYINPUT84), .ZN(n553) );
  NAND2_X1 U534 ( .A1(G902), .A2(n432), .ZN(n549) );
  NOR2_X1 U535 ( .A1(G900), .A2(n549), .ZN(n433) );
  AND2_X1 U536 ( .A1(n433), .A2(G953), .ZN(n434) );
  OR2_X1 U537 ( .A1(n553), .A2(n434), .ZN(n530) );
  INV_X1 U538 ( .A(n435), .ZN(n437) );
  INV_X1 U539 ( .A(G221), .ZN(n436) );
  OR2_X1 U540 ( .A1(n437), .A2(n436), .ZN(n439) );
  INV_X1 U541 ( .A(KEYINPUT21), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n599) );
  NAND2_X1 U543 ( .A1(n530), .A2(n599), .ZN(n440) );
  OR2_X1 U544 ( .A1(n600), .A2(n440), .ZN(n442) );
  INV_X1 U545 ( .A(KEYINPUT70), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n442), .B(n441), .ZN(n505) );
  NOR2_X1 U547 ( .A1(G953), .A2(G237), .ZN(n464) );
  NAND2_X1 U548 ( .A1(n464), .A2(G210), .ZN(n445) );
  XNOR2_X2 U549 ( .A(n443), .B(G143), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n494), .B(n734), .ZN(n481) );
  XNOR2_X1 U551 ( .A(G137), .B(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U552 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U553 ( .A(G902), .ZN(n489) );
  INV_X1 U554 ( .A(KEYINPUT72), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n450), .B(G472), .ZN(n451) );
  XNOR2_X1 U556 ( .A(n453), .B(KEYINPUT7), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n479), .B(n454), .ZN(n455) );
  XOR2_X1 U558 ( .A(n455), .B(KEYINPUT9), .Z(n460) );
  XNOR2_X1 U559 ( .A(n456), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U560 ( .A(n459), .B(n460), .ZN(n680) );
  NOR2_X1 U561 ( .A1(G902), .A2(n680), .ZN(n463) );
  XOR2_X1 U562 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n466) );
  NAND2_X1 U563 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U564 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U565 ( .A(G140), .B(G122), .Z(n468) );
  XNOR2_X1 U566 ( .A(G143), .B(G131), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n470), .B(n469), .ZN(n473) );
  XNOR2_X1 U569 ( .A(G113), .B(G104), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n477), .B(KEYINPUT12), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n670), .B(n471), .ZN(n472) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n561) );
  INV_X1 U574 ( .A(n561), .ZN(n503) );
  XNOR2_X1 U575 ( .A(n476), .B(G110), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n478), .B(n477), .ZN(n480) );
  NAND2_X1 U577 ( .A1(n725), .A2(G224), .ZN(n482) );
  XNOR2_X1 U578 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U580 ( .A(G237), .ZN(n488) );
  NAND2_X1 U581 ( .A1(n489), .A2(n488), .ZN(n493) );
  NAND2_X1 U582 ( .A1(n493), .A2(G210), .ZN(n491) );
  INV_X1 U583 ( .A(KEYINPUT78), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U585 ( .A1(n493), .A2(G214), .ZN(n611) );
  XNOR2_X1 U586 ( .A(n496), .B(n495), .ZN(n501) );
  NAND2_X1 U587 ( .A1(n725), .A2(G227), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n497), .B(G107), .ZN(n498) );
  XNOR2_X2 U589 ( .A(n502), .B(G469), .ZN(n511) );
  INV_X1 U590 ( .A(n555), .ZN(n575) );
  XNOR2_X1 U591 ( .A(n596), .B(KEYINPUT83), .ZN(n572) );
  NOR2_X1 U592 ( .A1(n719), .A2(n346), .ZN(n616) );
  INV_X1 U593 ( .A(n517), .ZN(n504) );
  NAND2_X1 U594 ( .A1(n505), .A2(n504), .ZN(n507) );
  XNOR2_X1 U595 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U597 ( .A1(n508), .A2(n511), .ZN(n528) );
  OR2_X1 U598 ( .A1(n528), .A2(n548), .ZN(n709) );
  NOR2_X1 U599 ( .A1(n616), .A2(n709), .ZN(n510) );
  XOR2_X1 U600 ( .A(KEYINPUT47), .B(n510), .Z(n523) );
  XNOR2_X1 U601 ( .A(n599), .B(KEYINPUT88), .ZN(n567) );
  AND2_X1 U602 ( .A1(n600), .A2(n567), .ZN(n597) );
  NAND2_X1 U603 ( .A1(n597), .A2(n511), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n512), .B(KEYINPUT89), .ZN(n579) );
  XNOR2_X1 U605 ( .A(n579), .B(KEYINPUT105), .ZN(n534) );
  INV_X1 U606 ( .A(n530), .ZN(n513) );
  NOR2_X1 U607 ( .A1(n561), .A2(n513), .ZN(n515) );
  NAND2_X1 U608 ( .A1(n515), .A2(n514), .ZN(n516) );
  NOR2_X1 U609 ( .A1(n562), .A2(n516), .ZN(n520) );
  INV_X1 U610 ( .A(n611), .ZN(n538) );
  OR2_X1 U611 ( .A1(n517), .A2(n538), .ZN(n519) );
  INV_X1 U612 ( .A(KEYINPUT30), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n519), .B(n518), .ZN(n532) );
  NAND2_X1 U614 ( .A1(n520), .A2(n532), .ZN(n521) );
  NOR2_X1 U615 ( .A1(n534), .A2(n521), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n522), .B(KEYINPUT106), .ZN(n653) );
  NOR2_X1 U617 ( .A1(n523), .A2(n653), .ZN(n524) );
  XNOR2_X1 U618 ( .A(n525), .B(KEYINPUT69), .ZN(n537) );
  XNOR2_X1 U619 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n514), .B(n526), .ZN(n612) );
  NAND2_X1 U621 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n614) );
  NOR2_X1 U623 ( .A1(n615), .A2(n614), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT41), .ZN(n630) );
  NOR2_X1 U625 ( .A1(n630), .A2(n528), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n529), .B(KEYINPUT42), .ZN(n740) );
  NAND2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U628 ( .A(n535), .B(KEYINPUT46), .ZN(n536) );
  NOR2_X1 U629 ( .A1(n596), .A2(n538), .ZN(n539) );
  AND2_X1 U630 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U631 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n541) );
  XNOR2_X1 U632 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U633 ( .A(KEYINPUT102), .B(n543), .ZN(n545) );
  INV_X1 U634 ( .A(n514), .ZN(n544) );
  NAND2_X1 U635 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U636 ( .A(n546), .B(KEYINPUT104), .ZN(n741) );
  NAND2_X1 U637 ( .A1(n547), .A2(n719), .ZN(n654) );
  INV_X1 U638 ( .A(n549), .ZN(n551) );
  INV_X1 U639 ( .A(G898), .ZN(n550) );
  AND2_X1 U640 ( .A1(n550), .A2(G953), .ZN(n736) );
  AND2_X1 U641 ( .A1(n551), .A2(n736), .ZN(n552) );
  OR2_X1 U642 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U643 ( .A1(n597), .A2(n555), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT99), .ZN(n556) );
  NAND2_X1 U645 ( .A1(n556), .A2(n571), .ZN(n558) );
  XNOR2_X1 U646 ( .A(KEYINPUT82), .B(KEYINPUT33), .ZN(n557) );
  XNOR2_X1 U647 ( .A(n558), .B(n557), .ZN(n620) );
  XNOR2_X1 U648 ( .A(n560), .B(n559), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U650 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U651 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n565) );
  INV_X1 U652 ( .A(n614), .ZN(n568) );
  XNOR2_X1 U653 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n569) );
  NOR2_X1 U654 ( .A1(n572), .A2(n600), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n588), .A2(n573), .ZN(n574) );
  XNOR2_X1 U656 ( .A(n576), .B(KEYINPUT64), .ZN(n577) );
  INV_X1 U657 ( .A(n600), .ZN(n586) );
  NOR2_X1 U658 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n578) );
  XNOR2_X1 U659 ( .A(n580), .B(KEYINPUT90), .ZN(n705) );
  OR2_X1 U660 ( .A1(n581), .A2(n517), .ZN(n582) );
  XNOR2_X1 U661 ( .A(n582), .B(KEYINPUT91), .ZN(n607) );
  XNOR2_X1 U662 ( .A(KEYINPUT92), .B(KEYINPUT31), .ZN(n583) );
  XNOR2_X1 U663 ( .A(n584), .B(n583), .ZN(n718) );
  NOR2_X1 U664 ( .A1(n705), .A2(n718), .ZN(n585) );
  NOR2_X1 U665 ( .A1(n585), .A2(n616), .ZN(n591) );
  NOR2_X1 U666 ( .A1(n586), .A2(n596), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n699) );
  NAND2_X1 U668 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n699), .A2(n589), .ZN(n590) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT50), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT49), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n517), .A2(n602), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT116), .ZN(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n630), .A2(n610), .ZN(n623) );
  NOR2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n618) );
  NOR2_X1 U683 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U684 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U685 ( .A(n619), .B(KEYINPUT118), .ZN(n621) );
  INV_X1 U686 ( .A(n620), .ZN(n629) );
  NOR2_X1 U687 ( .A1(n621), .A2(n629), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n623), .A2(n622), .ZN(n626) );
  NOR2_X1 U689 ( .A1(n628), .A2(n627), .ZN(n633) );
  NOR2_X1 U690 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U691 ( .A(n631), .B(KEYINPUT120), .ZN(n632) );
  NOR2_X1 U692 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U693 ( .A1(n640), .A2(n634), .ZN(n635) );
  NOR2_X1 U694 ( .A1(G953), .A2(n635), .ZN(n638) );
  XNOR2_X1 U695 ( .A(n636), .B(KEYINPUT53), .ZN(n637) );
  XNOR2_X1 U696 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n642) );
  XNOR2_X1 U697 ( .A(n642), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U698 ( .A(n641), .B(n643), .ZN(n644) );
  XNOR2_X1 U699 ( .A(n645), .B(n644), .ZN(n647) );
  INV_X1 U700 ( .A(G952), .ZN(n646) );
  NAND2_X1 U701 ( .A1(n646), .A2(G953), .ZN(n687) );
  NAND2_X1 U702 ( .A1(n692), .A2(G217), .ZN(n650) );
  XNOR2_X1 U703 ( .A(n648), .B(KEYINPUT125), .ZN(n649) );
  XNOR2_X1 U704 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U705 ( .A(G143), .B(n653), .Z(G45) );
  XNOR2_X1 U706 ( .A(n654), .B(G134), .ZN(G36) );
  XNOR2_X1 U707 ( .A(n655), .B(G110), .ZN(G12) );
  XOR2_X1 U708 ( .A(n656), .B(G119), .Z(G21) );
  XOR2_X1 U709 ( .A(G131), .B(n657), .Z(G33) );
  XOR2_X1 U710 ( .A(G125), .B(KEYINPUT37), .Z(n659) );
  XOR2_X1 U711 ( .A(n659), .B(n658), .Z(G27) );
  XOR2_X1 U712 ( .A(n660), .B(G122), .Z(G24) );
  NAND2_X1 U713 ( .A1(n692), .A2(G472), .ZN(n664) );
  XNOR2_X1 U714 ( .A(KEYINPUT108), .B(KEYINPUT62), .ZN(n661) );
  XNOR2_X1 U715 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U716 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U717 ( .A1(n665), .A2(n687), .ZN(n667) );
  XOR2_X1 U718 ( .A(KEYINPUT109), .B(KEYINPUT63), .Z(n666) );
  XNOR2_X1 U719 ( .A(n667), .B(n666), .ZN(G57) );
  INV_X1 U720 ( .A(n668), .ZN(n669) );
  XNOR2_X1 U721 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U722 ( .A(n672), .B(n671), .ZN(n675) );
  XOR2_X1 U723 ( .A(n675), .B(n673), .Z(n674) );
  NAND2_X1 U724 ( .A1(n674), .A2(n725), .ZN(n679) );
  XNOR2_X1 U725 ( .A(G227), .B(n675), .ZN(n676) );
  NAND2_X1 U726 ( .A1(n676), .A2(G900), .ZN(n677) );
  NAND2_X1 U727 ( .A1(G953), .A2(n677), .ZN(n678) );
  NAND2_X1 U728 ( .A1(n679), .A2(n678), .ZN(G72) );
  NAND2_X1 U729 ( .A1(n692), .A2(G478), .ZN(n682) );
  XNOR2_X1 U730 ( .A(n680), .B(KEYINPUT124), .ZN(n681) );
  XNOR2_X1 U731 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U732 ( .A(n687), .ZN(n697) );
  NOR2_X1 U733 ( .A1(n683), .A2(n697), .ZN(G63) );
  NAND2_X1 U734 ( .A1(n692), .A2(G475), .ZN(n686) );
  XOR2_X1 U735 ( .A(n684), .B(KEYINPUT59), .Z(n685) );
  XNOR2_X1 U736 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U737 ( .A1(n688), .A2(n687), .ZN(n691) );
  XNOR2_X1 U738 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n689) );
  XNOR2_X1 U739 ( .A(n689), .B(KEYINPUT66), .ZN(n690) );
  XNOR2_X1 U740 ( .A(n691), .B(n690), .ZN(G60) );
  NAND2_X1 U741 ( .A1(n692), .A2(G469), .ZN(n696) );
  XOR2_X1 U742 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U743 ( .A(n693), .B(n694), .ZN(n695) );
  XNOR2_X1 U744 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U745 ( .A1(n698), .A2(n697), .ZN(G54) );
  XNOR2_X1 U746 ( .A(G101), .B(n699), .ZN(G3) );
  NAND2_X1 U747 ( .A1(n705), .A2(n715), .ZN(n700) );
  XNOR2_X1 U748 ( .A(n700), .B(KEYINPUT110), .ZN(n701) );
  XNOR2_X1 U749 ( .A(G104), .B(n701), .ZN(G6) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n703) );
  XNOR2_X1 U751 ( .A(G107), .B(KEYINPUT26), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(n704) );
  XOR2_X1 U753 ( .A(KEYINPUT111), .B(n704), .Z(n707) );
  NAND2_X1 U754 ( .A1(n719), .A2(n705), .ZN(n706) );
  XNOR2_X1 U755 ( .A(n707), .B(n706), .ZN(G9) );
  XOR2_X1 U756 ( .A(n708), .B(KEYINPUT29), .Z(n711) );
  INV_X1 U757 ( .A(n709), .ZN(n712) );
  NAND2_X1 U758 ( .A1(n712), .A2(n719), .ZN(n710) );
  XNOR2_X1 U759 ( .A(n711), .B(n710), .ZN(G30) );
  XOR2_X1 U760 ( .A(G146), .B(KEYINPUT113), .Z(n714) );
  NAND2_X1 U761 ( .A1(n715), .A2(n712), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n714), .B(n713), .ZN(G48) );
  NAND2_X1 U763 ( .A1(n718), .A2(n715), .ZN(n716) );
  XNOR2_X1 U764 ( .A(n716), .B(KEYINPUT114), .ZN(n717) );
  XNOR2_X1 U765 ( .A(G113), .B(n717), .ZN(G15) );
  XOR2_X1 U766 ( .A(G116), .B(KEYINPUT115), .Z(n721) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n721), .B(n720), .ZN(G18) );
  INV_X1 U769 ( .A(n722), .ZN(n724) );
  NAND2_X1 U770 ( .A1(G898), .A2(KEYINPUT61), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U773 ( .A1(G224), .A2(KEYINPUT61), .ZN(n730) );
  AND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n727) );
  NOR2_X1 U775 ( .A1(KEYINPUT61), .A2(n727), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n550), .A2(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(KEYINPUT127), .ZN(n739) );
  XNOR2_X1 U780 ( .A(n734), .B(G101), .ZN(n735) );
  NOR2_X1 U781 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U782 ( .A(n739), .B(n738), .Z(G69) );
  XOR2_X1 U783 ( .A(G137), .B(n740), .Z(G39) );
  XNOR2_X1 U784 ( .A(G140), .B(n741), .ZN(G42) );
endmodule

