//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  AND2_X1   g0040(.A1(G1), .A2(G13), .ZN(new_n241));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n245));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n246), .B(G45), .C1(new_n244), .C2(KEYINPUT5), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n245), .B1(new_n247), .B2(KEYINPUT77), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT77), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT5), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G41), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n249), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(G270), .B(new_n243), .C1(new_n248), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT78), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n247), .A2(KEYINPUT77), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n251), .A2(new_n249), .A3(new_n253), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n241), .B2(new_n242), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n257), .A2(new_n258), .A3(new_n245), .A4(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n245), .A3(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT78), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n262), .A2(new_n263), .A3(G270), .A4(new_n243), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n256), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT65), .A3(new_n212), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT65), .B1(new_n266), .B2(new_n212), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n246), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G116), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G283), .ZN(new_n276));
  INV_X1    g0076(.A(G97), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n276), .B(new_n213), .C1(G33), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n266), .A2(new_n212), .ZN(new_n279));
  INV_X1    g0079(.A(G116), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT20), .A4(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(new_n271), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n284), .A2(new_n285), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G179), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  OAI211_X1 g0091(.A(G264), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  OAI211_X1 g0093(.A(G257), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(G303), .ZN(new_n295));
  OR2_X1    g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n243), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n265), .A2(new_n288), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n275), .B2(new_n287), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n300), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n256), .A2(new_n305), .A3(new_n261), .A4(new_n264), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT21), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n304), .B2(new_n306), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n306), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n311), .A2(new_n313), .A3(new_n288), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n298), .A2(G222), .A3(new_n293), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n298), .A2(G223), .A3(G1698), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n290), .A2(new_n291), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G77), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT64), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n243), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n321), .B2(new_n320), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n244), .A2(new_n250), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n246), .A2(new_n324), .B1(new_n241), .B2(new_n242), .ZN(new_n325));
  AOI21_X1  g0125(.A(G1), .B1(new_n244), .B2(new_n250), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(G226), .B1(new_n260), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n271), .A2(G50), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G20), .A2(G33), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT66), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n213), .A2(G33), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n330), .B1(new_n342), .B2(new_n270), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT65), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n279), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n267), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n246), .A2(G20), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G50), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n323), .A2(G190), .A3(new_n327), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n343), .A2(KEYINPUT9), .A3(new_n349), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n329), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT10), .ZN(new_n356));
  INV_X1    g0156(.A(new_n328), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n289), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n350), .C1(G169), .C2(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n226), .A2(G1698), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n360), .B1(G226), .B2(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G33), .A3(G97), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n300), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n260), .A2(new_n326), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n243), .A2(G238), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n243), .B1(new_n361), .B2(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n372), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT13), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G169), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n377), .A2(new_n383), .A3(new_n378), .A4(G169), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(G179), .A3(new_n376), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n380), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n346), .A2(new_n347), .ZN(new_n387));
  INV_X1    g0187(.A(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n271), .A2(G68), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT12), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n387), .A2(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(G20), .ZN(new_n394));
  INV_X1    g0194(.A(G77), .ZN(new_n395));
  INV_X1    g0195(.A(new_n331), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n394), .B1(new_n341), .B2(new_n395), .C1(new_n396), .C2(new_n202), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n270), .A2(new_n397), .A3(KEYINPUT11), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT11), .B1(new_n270), .B2(new_n397), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n393), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n373), .B2(new_n376), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n373), .A2(G190), .A3(new_n376), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n400), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n406), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT72), .B1(new_n408), .B2(new_n403), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n386), .A2(new_n401), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT8), .B(G58), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n411), .A2(new_n396), .B1(new_n213), .B2(new_n395), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n341), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n270), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n346), .A2(G77), .A3(new_n347), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n286), .A2(new_n395), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT69), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(G232), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT68), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n298), .A2(G238), .A3(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n318), .A2(G107), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n243), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n325), .A2(G244), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n370), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n303), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n424), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n423), .A2(new_n424), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n289), .B(new_n434), .C1(new_n437), .C2(new_n243), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n422), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n420), .A2(KEYINPUT70), .A3(new_n421), .ZN(new_n441));
  OAI21_X1  g0241(.A(G200), .B1(new_n430), .B2(new_n432), .ZN(new_n442));
  OAI211_X1 g0242(.A(G190), .B(new_n434), .C1(new_n437), .C2(new_n243), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT70), .B1(new_n420), .B2(new_n421), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n440), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n356), .A2(new_n359), .A3(new_n410), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n339), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n338), .A2(new_n335), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n271), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n348), .B2(new_n340), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT7), .B1(new_n318), .B2(new_n213), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n297), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(G68), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n334), .A2(new_n388), .ZN(new_n458));
  OAI21_X1  g0258(.A(G20), .B1(new_n458), .B2(new_n201), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n331), .A2(G159), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n453), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n296), .A2(new_n213), .A3(new_n297), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT7), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n388), .B1(new_n466), .B2(new_n455), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(KEYINPUT16), .A3(new_n460), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n270), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n452), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G223), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n293), .ZN(new_n472));
  INV_X1    g0272(.A(G226), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n474), .C1(new_n290), .C2(new_n291), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n300), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n325), .A2(G232), .B1(new_n260), .B2(new_n326), .ZN(new_n479));
  AOI21_X1  g0279(.A(G169), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT75), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n477), .B2(new_n300), .ZN(new_n482));
  AOI211_X1 g0282(.A(KEYINPUT75), .B(new_n243), .C1(new_n475), .C2(new_n476), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n243), .A2(G232), .A3(new_n371), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n370), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G179), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n480), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n470), .A2(new_n488), .A3(KEYINPUT18), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT76), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT76), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n470), .A2(new_n488), .A3(new_n491), .A4(KEYINPUT18), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT18), .ZN(new_n493));
  INV_X1    g0293(.A(new_n468), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n346), .B1(new_n457), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n453), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n467), .B2(new_n461), .ZN(new_n497));
  INV_X1    g0297(.A(new_n340), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n387), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n497), .B1(new_n499), .B2(new_n451), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n243), .B1(new_n475), .B2(new_n476), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n481), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n487), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n480), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n493), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n490), .A2(new_n492), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n486), .A2(G190), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n501), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  AOI21_X1  g0310(.A(G200), .B1(new_n478), .B2(new_n479), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n500), .A2(new_n513), .A3(KEYINPUT17), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT17), .B1(new_n500), .B2(new_n513), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n448), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n520));
  OAI211_X1 g0320(.A(G238), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n521));
  INV_X1    g0321(.A(G33), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n280), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n525), .A2(new_n300), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n246), .A2(new_n259), .A3(G45), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n250), .B2(G1), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n243), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n303), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n525), .B2(new_n300), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n289), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n413), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n274), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n271), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  INV_X1    g0340(.A(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n277), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n363), .B2(new_n365), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n544), .B2(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n296), .B2(new_n297), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(G68), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n537), .B(new_n539), .C1(new_n549), .C2(new_n346), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n533), .A2(new_n402), .ZN(new_n551));
  AOI211_X1 g0351(.A(new_n312), .B(new_n531), .C1(new_n525), .C2(new_n300), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n346), .B1(new_n545), .B2(new_n548), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n270), .A2(new_n540), .A3(new_n273), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n554), .A2(new_n555), .A3(new_n538), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n535), .A2(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n298), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n298), .A2(G250), .A3(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n276), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n300), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n262), .A2(G257), .A3(new_n243), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n261), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n567), .A2(new_n277), .A3(G107), .ZN(new_n568));
  XNOR2_X1  g0368(.A(G97), .B(G107), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(new_n213), .B1(new_n395), .B2(new_n396), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n541), .B1(new_n466), .B2(new_n455), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n270), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n273), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n346), .A2(G97), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n286), .A2(new_n277), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n566), .A2(new_n303), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n564), .A2(new_n289), .A3(new_n261), .A4(new_n565), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n575), .B1(G97), .B2(new_n271), .ZN(new_n581));
  INV_X1    g0381(.A(new_n572), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n569), .A2(new_n567), .ZN(new_n583));
  INV_X1    g0383(.A(new_n568), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(G20), .B1(G77), .B2(new_n331), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n581), .B1(new_n587), .B2(new_n270), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n564), .A2(G190), .A3(new_n261), .A4(new_n565), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n564), .A2(new_n261), .A3(new_n565), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n402), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n557), .A2(new_n580), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n213), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n541), .A2(KEYINPUT23), .A3(G20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n523), .A2(new_n213), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n546), .A2(G87), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n213), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n601));
  XOR2_X1   g0401(.A(KEYINPUT79), .B(KEYINPUT22), .Z(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n598), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n270), .B1(new_n604), .B2(KEYINPUT24), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n606), .B(new_n598), .C1(new_n600), .C2(new_n603), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n574), .B(G107), .C1(new_n268), .C2(new_n269), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT80), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n246), .A2(new_n541), .A3(G13), .A4(G20), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT25), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n608), .B2(new_n612), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n605), .A2(new_n607), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n616));
  OAI211_X1 g0416(.A(G250), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G294), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n300), .ZN(new_n620));
  OAI211_X1 g0420(.A(G264), .B(new_n243), .C1(new_n248), .C2(new_n254), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n261), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(G179), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n303), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n402), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n620), .A2(new_n621), .A3(new_n312), .A4(new_n261), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n613), .A2(new_n614), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n600), .A2(new_n603), .ZN(new_n630));
  INV_X1    g0430(.A(new_n598), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n606), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n604), .A2(KEYINPUT24), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n270), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n629), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT81), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n625), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n625), .B2(new_n636), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n315), .A2(new_n519), .A3(new_n592), .A4(new_n640), .ZN(G372));
  NAND3_X1  g0441(.A1(new_n550), .A2(new_n532), .A3(new_n534), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n557), .A2(new_n580), .A3(new_n591), .A4(new_n636), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n625), .B(new_n302), .C1(new_n308), .C2(new_n309), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n553), .A2(new_n556), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(new_n578), .A3(new_n642), .A4(new_n579), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT82), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n578), .A2(new_n579), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT82), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n557), .A3(new_n652), .A4(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n649), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n519), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n359), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n507), .A2(new_n489), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n409), .A2(new_n407), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n440), .B1(new_n386), .B2(new_n401), .ZN(new_n661));
  INV_X1    g0461(.A(new_n516), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n514), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n664), .B2(new_n356), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(G369));
  NAND3_X1  g0466(.A1(new_n246), .A2(new_n213), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n615), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n625), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n288), .A2(new_n672), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n315), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n310), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n672), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n640), .A2(new_n310), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n672), .B(KEYINPUT83), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n675), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  NOR2_X1   g0491(.A1(new_n542), .A2(G116), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n207), .A2(new_n244), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(G1), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n210), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n648), .B(new_n649), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n672), .B1(new_n646), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(new_n688), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n646), .B2(new_n655), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(KEYINPUT29), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n640), .A2(new_n315), .A3(new_n592), .A4(new_n688), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n533), .A2(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n566), .A2(new_n306), .A3(new_n622), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n301), .A2(new_n533), .A3(new_n621), .A4(new_n620), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n256), .A2(new_n261), .A3(new_n264), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n566), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(KEYINPUT30), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT85), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n711), .A3(KEYINPUT30), .ZN(new_n712));
  AND4_X1   g0512(.A1(new_n301), .A2(new_n533), .A3(new_n621), .A4(new_n620), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n590), .A2(new_n713), .A3(new_n265), .A4(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT85), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n704), .B1(new_n716), .B2(new_n686), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n710), .A2(KEYINPUT84), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n715), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT84), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(new_n706), .C1(new_n709), .C2(KEYINPUT30), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n688), .A2(new_n704), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n703), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n702), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(new_n683), .ZN(new_n730));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n246), .B1(new_n732), .B2(G45), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(new_n693), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT86), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n682), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n298), .A2(new_n207), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n739), .B1(G116), .B2(new_n207), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n236), .A2(new_n250), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n318), .A2(new_n207), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n250), .B2(new_n211), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT87), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n212), .B1(G20), .B2(new_n303), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n213), .A2(new_n289), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n312), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n213), .A2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n289), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n298), .B1(new_n762), .B2(G311), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n764), .B1(G326), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n289), .A2(new_n402), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT89), .ZN(new_n769));
  OAI21_X1  g0569(.A(G20), .B1(new_n769), .B2(new_n312), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G294), .ZN(new_n771));
  INV_X1    g0571(.A(new_n759), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n213), .A2(new_n312), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n402), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n760), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n295), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n759), .A2(new_n776), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G283), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n767), .A2(new_n771), .A3(new_n774), .A4(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n753), .A2(new_n388), .B1(new_n765), .B2(new_n202), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n395), .A2(new_n761), .B1(new_n781), .B2(new_n541), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n298), .B1(new_n777), .B2(new_n540), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n778), .B(KEYINPUT88), .Z(new_n789));
  INV_X1    g0589(.A(new_n770), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n789), .B2(new_n334), .C1(new_n790), .C2(new_n277), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n773), .A2(G159), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n784), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n751), .B1(new_n794), .B2(new_n748), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  INV_X1    g0596(.A(new_n747), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n682), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n737), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  INV_X1    g0600(.A(KEYINPUT70), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n422), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n802), .A2(new_n441), .A3(new_n443), .A4(new_n442), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n422), .A2(new_n672), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n440), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n439), .A2(new_n672), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n805), .A2(new_n700), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n808));
  INV_X1    g0608(.A(new_n645), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n557), .A2(new_n580), .A3(new_n591), .A4(new_n636), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n642), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n807), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n806), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n446), .A2(new_n441), .B1(new_n422), .B2(new_n672), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n440), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n812), .B1(new_n701), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n735), .B1(new_n817), .B2(new_n726), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n726), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(new_n748), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n766), .A2(G137), .B1(new_n762), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n753), .ZN(new_n823));
  INV_X1    g0623(.A(new_n789), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(G143), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT34), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n298), .B1(new_n781), .B2(new_n388), .C1(new_n202), .C2(new_n777), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G132), .B2(new_n773), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n334), .B2(new_n790), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n765), .A2(new_n295), .B1(new_n761), .B2(new_n280), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G283), .B2(new_n754), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT92), .Z(new_n832));
  OAI21_X1  g0632(.A(new_n318), .B1(new_n777), .B2(new_n541), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT93), .Z(new_n834));
  AOI22_X1  g0634(.A1(new_n773), .A2(G311), .B1(G87), .B2(new_n782), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n778), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n770), .A2(G97), .B1(G294), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT94), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n826), .A2(new_n829), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n820), .B1(new_n840), .B2(KEYINPUT95), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(KEYINPUT95), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n735), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n748), .A2(new_n745), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT91), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n843), .B1(new_n395), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n842), .B(new_n847), .C1(new_n746), .C2(new_n816), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n819), .A2(new_n848), .ZN(G384));
  OR2_X1    g0649(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n214), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI211_X1 g0653(.A(new_n211), .B(G77), .C1(new_n334), .C2(new_n388), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n246), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n386), .A2(new_n401), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n672), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n500), .A2(new_n670), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n508), .B2(new_n517), .ZN(new_n864));
  NOR2_X1   g0664(.A1(KEYINPUT97), .A2(KEYINPUT37), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n511), .B1(new_n484), .B2(new_n509), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT97), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n470), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n495), .A2(new_n497), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n506), .A2(new_n670), .B1(new_n870), .B2(new_n452), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n865), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n500), .A2(new_n513), .B1(KEYINPUT97), .B2(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(new_n670), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n470), .B1(new_n488), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n865), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n861), .B1(new_n864), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n518), .A2(new_n862), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT98), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT98), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n864), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n880), .A2(new_n882), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n863), .B1(new_n517), .B2(new_n659), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n861), .B1(new_n889), .B2(new_n878), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n860), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n409), .A2(new_n407), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n401), .B(new_n672), .C1(new_n894), .C2(new_n386), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n401), .A2(new_n672), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n858), .A2(new_n660), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n688), .B(new_n813), .C1(new_n814), .C2(new_n440), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n646), .B2(new_n655), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n806), .B(KEYINPUT96), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n869), .A2(new_n871), .A3(new_n865), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n876), .B1(new_n873), .B2(new_n875), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n880), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n884), .B1(new_n864), .B2(new_n881), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT98), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n902), .A2(new_n909), .B1(new_n659), .B2(new_n874), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT99), .B1(new_n893), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n895), .A2(new_n897), .ZN(new_n912));
  INV_X1    g0712(.A(new_n901), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n812), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n659), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n886), .B1(new_n915), .B2(new_n670), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT99), .ZN(new_n917));
  INV_X1    g0717(.A(new_n892), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(KEYINPUT39), .B2(new_n886), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n916), .B(new_n917), .C1(new_n919), .C2(new_n860), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n519), .B(new_n699), .C1(KEYINPUT29), .C2(new_n701), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n665), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT100), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n712), .A2(new_n715), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT31), .B(new_n672), .C1(new_n926), .C2(new_n710), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n703), .A2(new_n717), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n815), .B1(new_n895), .B2(new_n897), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n862), .B1(new_n915), .B2(new_n663), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n931), .B2(new_n905), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n864), .A2(new_n881), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT40), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n925), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n888), .B2(new_n890), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n937), .A2(KEYINPUT100), .A3(new_n928), .A4(new_n929), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n886), .A2(new_n928), .A3(new_n929), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n935), .A2(new_n938), .B1(new_n939), .B2(new_n936), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n519), .A2(new_n928), .ZN(new_n942));
  OAI21_X1  g0742(.A(G330), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n924), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(G1), .B1(new_n731), .B2(G20), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(KEYINPUT101), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n944), .B2(new_n924), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT101), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n857), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NOR2_X1   g0750(.A1(new_n556), .A2(new_n686), .ZN(new_n951));
  MUX2_X1   g0751(.A(new_n557), .B(new_n643), .S(new_n951), .Z(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n580), .B(new_n591), .C1(new_n588), .C2(new_n688), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n651), .A2(new_n700), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n687), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n580), .B1(new_n954), .B2(new_n625), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(KEYINPUT42), .B1(new_n688), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n953), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n952), .A2(KEYINPUT102), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n952), .A2(KEYINPUT102), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT104), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n962), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n968), .B1(new_n962), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n685), .A2(new_n957), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n970), .B2(new_n971), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n693), .B(KEYINPUT41), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT105), .B1(new_n690), .B2(new_n956), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n687), .A2(new_n689), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT105), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n957), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n978), .A2(new_n957), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT45), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n980), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n684), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n983), .A2(new_n985), .A3(new_n685), .A4(new_n986), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n674), .B(new_n676), .C1(new_n681), .C2(new_n672), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n683), .A2(new_n990), .A3(new_n687), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n683), .B1(new_n990), .B2(new_n687), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n727), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n976), .B1(new_n995), .B2(new_n728), .ZN(new_n996));
  INV_X1    g0796(.A(new_n733), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n975), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n749), .B1(new_n207), .B2(new_n413), .C1(new_n232), .C2(new_n742), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n735), .ZN(new_n1000));
  INV_X1    g0800(.A(G159), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n298), .B1(new_n777), .B2(new_n334), .C1(new_n1001), .C2(new_n753), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n766), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n770), .A2(G68), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT106), .B(G137), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n773), .A2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n778), .A2(new_n822), .B1(new_n761), .B2(new_n202), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G77), .B2(new_n782), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n777), .A2(new_n280), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT46), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G311), .B2(new_n766), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(KEYINPUT46), .A2(new_n1010), .B1(new_n754), .B2(G294), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n541), .C2(new_n790), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n781), .A2(new_n277), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n298), .B(new_n1015), .C1(G283), .C2(new_n762), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n773), .A2(G317), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n295), .C2(new_n789), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1009), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n1000), .B1(new_n952), .B2(new_n797), .C1(new_n1020), .C2(new_n820), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n998), .A2(new_n1021), .ZN(G387));
  XNOR2_X1  g0822(.A(new_n693), .B(KEYINPUT112), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n994), .A2(KEYINPUT113), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n993), .A2(new_n727), .ZN(new_n1026));
  OAI21_X1  g0826(.A(KEYINPUT113), .B1(new_n994), .B2(new_n1024), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n993), .A2(KEYINPUT107), .A3(new_n733), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT107), .B1(new_n993), .B2(new_n733), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n678), .A2(new_n747), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n754), .A2(G311), .B1(new_n762), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n779), .B2(new_n765), .C1(new_n789), .C2(new_n755), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n777), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n770), .A2(G283), .B1(G294), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n318), .B1(new_n781), .B2(new_n280), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n773), .B2(G326), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n770), .A2(new_n536), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n202), .B2(new_n778), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT110), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n340), .A2(new_n753), .B1(new_n388), .B2(new_n761), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT111), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n318), .B(new_n1015), .C1(G77), .C2(new_n1037), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1001), .B2(new_n765), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G150), .B2(new_n773), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n820), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n229), .A2(G45), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT108), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n692), .ZN(new_n1058));
  AOI211_X1 g0858(.A(G45), .B(new_n1058), .C1(G68), .C2(G77), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n411), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n742), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(G107), .B2(new_n207), .C1(new_n692), .C2(new_n738), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n843), .B(new_n1055), .C1(new_n749), .C2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1028), .A2(new_n1067), .ZN(G393));
  NAND3_X1  g0868(.A1(new_n988), .A2(new_n997), .A3(new_n989), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n749), .B1(new_n277), .B2(new_n207), .C1(new_n239), .C2(new_n742), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n735), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n765), .A2(new_n822), .B1(new_n778), .B2(new_n1001), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT114), .Z(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n777), .A2(new_n388), .B1(new_n761), .B2(new_n411), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n318), .B(new_n1075), .C1(G87), .C2(new_n782), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n770), .A2(G77), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n773), .A2(G143), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n754), .A2(G50), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n773), .A2(G322), .B1(G283), .B2(new_n1037), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT116), .Z(new_n1082));
  AOI22_X1  g0882(.A1(new_n766), .A2(G317), .B1(new_n837), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(G294), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n318), .B1(new_n761), .B2(new_n1086), .C1(new_n541), .C2(new_n781), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G303), .B2(new_n754), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(new_n280), .C2(new_n790), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1074), .A2(new_n1080), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1071), .B1(new_n1090), .B2(new_n748), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n956), .B2(new_n797), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n995), .A2(new_n1023), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n994), .B1(new_n988), .B2(new_n989), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1069), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(G390));
  AND2_X1   g0895(.A1(new_n928), .A2(G330), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n519), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n922), .A3(new_n665), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n812), .A2(new_n913), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n725), .A2(G330), .A3(new_n816), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n912), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n928), .A2(new_n929), .A3(G330), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n928), .A2(G330), .A3(new_n816), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n912), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n901), .B1(new_n698), .B2(new_n816), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n725), .A2(G330), .A3(new_n816), .A4(new_n898), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1098), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n859), .B1(new_n888), .B2(new_n890), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1106), .B2(new_n912), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n892), .B1(new_n909), .B2(new_n891), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n859), .B1(new_n1099), .B2(new_n898), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1102), .A2(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1107), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n928), .A2(new_n929), .A3(new_n1119), .A4(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1110), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1097), .A2(new_n922), .A3(new_n665), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1096), .A2(new_n929), .B1(new_n1100), .B2(new_n912), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1099), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1108), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1117), .A2(new_n1122), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1023), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1123), .A2(new_n733), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n735), .B1(new_n845), .B2(new_n498), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1113), .A2(new_n746), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n318), .B1(new_n777), .B2(new_n540), .C1(new_n541), .C2(new_n753), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G283), .B2(new_n766), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n773), .A2(G294), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n388), .A2(new_n781), .B1(new_n761), .B2(new_n277), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G116), .B2(new_n837), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1077), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1037), .A2(G150), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT53), .Z(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n765), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n754), .B2(new_n1005), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n773), .A2(G125), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n781), .A2(new_n202), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n298), .B1(new_n761), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G132), .C2(new_n837), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n790), .A2(new_n1001), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1139), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT118), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n820), .B1(new_n1152), .B2(KEYINPUT118), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1132), .B(new_n1133), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1131), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1130), .A2(new_n1156), .ZN(G378));
  NOR2_X1   g0957(.A1(G33), .A2(G41), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT119), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G50), .B(new_n1159), .C1(new_n244), .C2(new_n318), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G41), .B(new_n298), .C1(new_n1037), .C2(G77), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n277), .B2(new_n753), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G116), .B2(new_n766), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n536), .A2(new_n762), .B1(new_n782), .B2(G58), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n541), .B2(new_n778), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G283), .B2(new_n773), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1004), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1142), .A2(new_n778), .B1(new_n777), .B2(new_n1147), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G137), .B2(new_n762), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n754), .A2(G132), .B1(new_n766), .B2(G125), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n790), .C2(new_n822), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1159), .B1(new_n1001), .B2(new_n781), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n773), .B2(G124), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1169), .B1(new_n1168), .B2(new_n1167), .C1(new_n1174), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n748), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n843), .B1(new_n202), .B2(new_n846), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n356), .A2(new_n359), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n350), .A2(new_n874), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  AND2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1183), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1182), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1180), .B(new_n1181), .C1(new_n1194), .C2(new_n746), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n940), .B2(G330), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n935), .A2(new_n938), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n936), .B1(new_n909), .B2(new_n930), .ZN(new_n1199));
  AND4_X1   g0999(.A1(G330), .A2(new_n1198), .A3(new_n1199), .A4(new_n1193), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n921), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(G330), .A3(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1194), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1198), .A2(new_n1193), .A3(G330), .A4(new_n1199), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1203), .A2(new_n920), .A3(new_n911), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1196), .B1(new_n1206), .B2(new_n997), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1201), .A2(new_n1205), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1023), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1129), .A2(new_n1125), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1209), .B2(new_n1211), .ZN(G375));
  NOR2_X1   g1012(.A1(new_n1128), .A2(new_n1125), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1213), .A2(new_n1109), .A3(new_n976), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT121), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n733), .B(KEYINPUT122), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n912), .A2(new_n745), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n735), .B1(new_n845), .B2(G68), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n318), .B1(new_n781), .B2(new_n395), .C1(new_n765), .C2(new_n1086), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G116), .B2(new_n754), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n773), .A2(G303), .ZN(new_n1221));
  INV_X1    g1021(.A(G283), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n778), .A2(new_n1222), .B1(new_n761), .B2(new_n541), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G97), .B2(new_n1037), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1046), .A3(new_n1221), .A4(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n824), .A2(new_n1005), .B1(G128), .B2(new_n773), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n777), .A2(new_n1001), .B1(new_n761), .B2(new_n822), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n318), .B(new_n1227), .C1(G58), .C2(new_n782), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n753), .C2(new_n1147), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n766), .A2(G132), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n202), .B2(new_n790), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1225), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1218), .B1(new_n1233), .B2(new_n748), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1128), .A2(new_n1216), .B1(new_n1217), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1215), .A2(new_n1235), .ZN(G381));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  INV_X1    g1037(.A(G390), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G387), .A2(new_n1241), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n671), .A2(G213), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1237), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G375), .C2(new_n1245), .ZN(G409));
  AOI21_X1  g1046(.A(new_n799), .B1(new_n1028), .B2(new_n1067), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1240), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n998), .A2(new_n1021), .A3(G390), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n998), .B2(new_n1021), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1238), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1240), .A2(new_n1247), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n998), .A2(new_n1021), .A3(G390), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G378), .B(new_n1207), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1206), .A2(new_n1216), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1195), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n976), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1206), .A2(new_n1260), .A3(new_n1210), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1237), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1128), .B2(new_n1125), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n1213), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1103), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1268));
  OAI211_X1 g1068(.A(KEYINPUT124), .B(new_n1268), .C1(new_n1109), .C2(new_n1265), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1024), .B1(new_n1213), .B2(KEYINPUT60), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1235), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1239), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1235), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1263), .A2(new_n1243), .A3(new_n1276), .ZN(new_n1277));
  XOR2_X1   g1077(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1278));
  AOI21_X1  g1078(.A(new_n1256), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1244), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1281), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1244), .A2(G2897), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1244), .A2(KEYINPUT126), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1273), .A2(new_n1274), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1273), .A2(new_n1274), .A3(new_n1285), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1286), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1280), .B1(new_n1292), .B2(new_n1281), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1294));
  AND4_X1   g1094(.A1(new_n1243), .A2(new_n1263), .A3(new_n1276), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1281), .B2(new_n1276), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1293), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1256), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1291), .B1(new_n1299), .B2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1237), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1275), .B1(new_n1302), .B2(new_n1257), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1275), .A3(new_n1257), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1256), .ZN(G402));
endmodule


