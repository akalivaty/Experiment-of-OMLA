//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n204), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(G50), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n209), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n216), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  INV_X1    g0037(.A(G107), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G97), .ZN(new_n239));
  INV_X1    g0039(.A(G97), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n220), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G20), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G50), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G50), .B2(new_n246), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT66), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n204), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G50), .A2(G58), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n204), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(G223), .B1(new_n273), .B2(G77), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n220), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  INV_X1    g0086(.A(new_n220), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n285), .A2(G226), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n280), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n266), .B1(new_n294), .B2(G169), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n293), .A2(G179), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n255), .A2(KEYINPUT9), .A3(new_n265), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT74), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n266), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n302), .A2(new_n303), .B1(new_n294), .B2(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n301), .A2(new_n306), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n299), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n257), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G77), .B1(G20), .B2(new_n263), .ZN(new_n314));
  INV_X1    g0114(.A(G50), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n260), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n247), .A2(new_n263), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n250), .A2(G68), .A3(new_n251), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT11), .B1(new_n316), .B2(new_n249), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(G232), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n325));
  OAI211_X1 g0125(.A(G226), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n279), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n285), .A2(G238), .B1(new_n288), .B2(new_n291), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(G179), .A3(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n329), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g0137(.A(G169), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n338), .B2(KEYINPUT14), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(new_n334), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n324), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G200), .B1(new_n336), .B2(new_n337), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n332), .A2(G190), .A3(new_n334), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n323), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT70), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n257), .ZN(new_n353));
  INV_X1    g0153(.A(G77), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n256), .A2(new_n260), .B1(new_n204), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n249), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  INV_X1    g0157(.A(new_n249), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n246), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n251), .A2(G77), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n250), .A2(KEYINPUT71), .A3(G77), .A4(new_n251), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n247), .A2(new_n354), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n356), .A2(KEYINPUT72), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n350), .B(KEYINPUT70), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n355), .B1(new_n366), .B2(new_n313), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n363), .B(new_n364), .C1(new_n367), .C2(new_n358), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n291), .A2(new_n282), .A3(G274), .ZN(new_n371));
  INV_X1    g0171(.A(G244), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n284), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(G238), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n268), .A2(new_n269), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n238), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT68), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n275), .A2(new_n378), .A3(G232), .ZN(new_n379));
  OAI211_X1 g0179(.A(G232), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT68), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT69), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n279), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n381), .ZN(new_n385));
  INV_X1    g0185(.A(new_n377), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(KEYINPUT69), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n374), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n365), .B(new_n370), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n282), .B1(new_n387), .B2(KEYINPUT69), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n382), .A2(new_n383), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n373), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n374), .C1(new_n384), .C2(new_n388), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n368), .C1(new_n394), .C2(G169), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n312), .A2(new_n349), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G1698), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(G223), .B2(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n279), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n285), .A2(G232), .B1(new_n288), .B2(new_n291), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n398), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G169), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n282), .B1(new_n406), .B2(new_n407), .ZN(new_n413));
  INV_X1    g0213(.A(G232), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n371), .B1(new_n414), .B2(new_n284), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n412), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n268), .A2(new_n204), .A3(new_n269), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n263), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G58), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n263), .ZN(new_n425));
  OAI21_X1  g0225(.A(G20), .B1(new_n425), .B2(new_n218), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n259), .A2(G159), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT7), .B1(new_n273), .B2(new_n204), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n271), .A2(new_n272), .A3(new_n420), .A4(G20), .ZN(new_n431));
  OAI21_X1  g0231(.A(G68), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n428), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(KEYINPUT16), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n434), .A3(new_n249), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n256), .B1(new_n203), .B2(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n250), .B1(new_n247), .B2(new_n256), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT18), .B(new_n417), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n437), .ZN(new_n440));
  INV_X1    g0240(.A(new_n417), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT75), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n437), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n432), .A2(new_n433), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n358), .B1(new_n445), .B2(new_n418), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(new_n434), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n447), .B2(new_n417), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n440), .A2(new_n439), .A3(new_n441), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n409), .A2(new_n390), .A3(new_n410), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n395), .B1(new_n413), .B2(new_n415), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n435), .A2(new_n437), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n435), .A2(KEYINPUT17), .A3(new_n454), .A4(new_n437), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n443), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n403), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n239), .A3(new_n241), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n239), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(KEYINPUT77), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n240), .A2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(new_n463), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(KEYINPUT77), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT78), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n470), .A4(new_n464), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(G20), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n238), .B1(new_n421), .B2(new_n422), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(G77), .B2(new_n259), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n249), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n246), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n203), .A2(G33), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n358), .A2(new_n246), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n372), .A2(G1698), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(KEYINPUT4), .C1(new_n272), .C2(new_n271), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n376), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G250), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n267), .A2(G244), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n268), .B2(new_n269), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n494), .B(new_n495), .C1(new_n497), .C2(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n279), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n290), .A2(G1), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT5), .B(G41), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n288), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G257), .A3(new_n282), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT80), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT80), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n499), .A2(new_n398), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT80), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT80), .B1(new_n502), .B2(new_n506), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .A3(new_n398), .A4(new_n499), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n499), .A2(new_n509), .A3(new_n510), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n412), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n487), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n499), .A2(new_n509), .A3(new_n510), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n482), .A3(new_n486), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n366), .A2(new_n485), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT83), .B(G87), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n204), .B1(new_n327), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n257), .B2(new_n240), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n376), .A2(new_n204), .A3(G68), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n249), .B1(new_n247), .B2(new_n352), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n288), .A2(new_n500), .ZN(new_n537));
  INV_X1    g0337(.A(G250), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n203), .B2(G45), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n282), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n539), .B2(new_n282), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g0344(.A1(G238), .A2(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n372), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n271), .C2(new_n272), .ZN(new_n547));
  INV_X1    g0347(.A(G33), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n282), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G169), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n282), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n541), .B1(new_n288), .B2(new_n500), .ZN(new_n556));
  INV_X1    g0356(.A(new_n552), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(G179), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n526), .A2(new_n536), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n557), .A3(G190), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT84), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n485), .A2(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n536), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n395), .B1(new_n556), .B2(new_n557), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n559), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n521), .A2(new_n525), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT85), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n521), .A2(KEYINPUT85), .A3(new_n525), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n204), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n238), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n550), .B2(new_n204), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n376), .A2(new_n204), .A3(G87), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n249), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n485), .A2(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT25), .B1(new_n247), .B2(new_n238), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT88), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n275), .A2(new_n591), .A3(G250), .ZN(new_n592));
  OAI211_X1 g0392(.A(G250), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT88), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G294), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n282), .B1(new_n600), .B2(KEYINPUT89), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n592), .B2(new_n594), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT89), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n279), .B1(new_n500), .B2(new_n501), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n601), .A2(new_n604), .B1(G264), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n398), .A3(new_n502), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(G264), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n279), .B1(new_n602), .B2(new_n603), .ZN(new_n609));
  AOI211_X1 g0409(.A(KEYINPUT89), .B(new_n598), .C1(new_n594), .C2(new_n592), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n502), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n412), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n590), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(G200), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n600), .A2(KEYINPUT89), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n604), .A3(new_n279), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(G190), .A3(new_n502), .A4(new_n608), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n584), .A4(new_n589), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n505), .A2(G270), .A3(new_n282), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT86), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT86), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n505), .A2(new_n622), .A3(G270), .A4(new_n282), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(G274), .B1(new_n278), .B2(new_n220), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n505), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G264), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n627));
  OAI211_X1 g0427(.A(G257), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n268), .A2(G303), .A3(new_n269), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n626), .B1(new_n630), .B2(new_n279), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT87), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n246), .B2(G116), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n247), .A2(KEYINPUT87), .A3(new_n549), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n485), .A2(G116), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n495), .B(new_n204), .C1(G33), .C2(new_n240), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n549), .A2(G20), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n249), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n632), .A2(G179), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n412), .B1(new_n636), .B2(new_n641), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT21), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n624), .A2(new_n631), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n632), .A2(new_n395), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n646), .A2(new_n390), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n642), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n461), .A2(new_n571), .A3(new_n619), .A4(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n559), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n564), .B(KEYINPUT90), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n536), .A2(new_n560), .A3(new_n562), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n559), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n618), .A2(new_n521), .A3(new_n525), .A4(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n584), .A2(new_n589), .B1(new_n611), .B2(new_n412), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n649), .B1(new_n660), .B2(new_n607), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n513), .A2(new_n517), .B1(new_n412), .B2(new_n519), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n566), .A2(new_n487), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n658), .A2(new_n666), .A3(new_n487), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n461), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n309), .A2(new_n311), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n438), .A2(new_n442), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n344), .B1(new_n347), .B2(new_n401), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n457), .A2(new_n458), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n299), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(KEYINPUT27), .B2(new_n678), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(G343), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n642), .ZN(new_n688));
  MUX2_X1   g0488(.A(new_n649), .B(new_n653), .S(new_n688), .Z(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n613), .A2(new_n618), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n584), .B2(new_n589), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n613), .B2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n649), .A2(new_n686), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n686), .B(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n613), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0503(.A(new_n207), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n529), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n219), .A2(G50), .A3(new_n222), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n669), .A2(new_n698), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n658), .A2(new_n487), .A3(new_n663), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT26), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(KEYINPUT26), .B2(new_n664), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n686), .C1(new_n718), .C2(new_n662), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n653), .A2(new_n613), .A3(new_n618), .A4(new_n698), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n571), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n544), .A2(new_n398), .A3(new_n552), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n632), .A2(new_n499), .A3(new_n516), .A4(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT30), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n519), .A2(new_n558), .A3(new_n646), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n606), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n556), .B2(new_n557), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT95), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n732), .A2(new_n646), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n732), .B2(new_n646), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n522), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n728), .A2(new_n731), .B1(new_n736), .B2(new_n611), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n724), .B1(new_n737), .B2(new_n686), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n699), .A2(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n731), .A2(new_n728), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n735), .A2(new_n522), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n732), .A2(new_n646), .A3(new_n733), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n611), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n738), .A2(new_n745), .A3(KEYINPUT96), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT96), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n730), .B1(new_n729), .B2(new_n606), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT30), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n750), .B2(new_n687), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n747), .B1(new_n751), .B2(new_n744), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n723), .A2(new_n746), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n720), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n712), .B1(new_n756), .B2(G1), .ZN(G364));
  AND2_X1   g0557(.A1(new_n204), .A2(G13), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n203), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n705), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n691), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n689), .ZN(new_n763));
  INV_X1    g0563(.A(new_n761), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n236), .A2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n704), .A2(new_n376), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n765), .B(new_n766), .C1(G45), .C2(new_n709), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n704), .A2(new_n273), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n768), .A2(G355), .B1(new_n549), .B2(new_n704), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n220), .B1(G20), .B2(new_n412), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n764), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  INV_X1    g0577(.A(new_n774), .ZN(new_n778));
  OAI21_X1  g0578(.A(G20), .B1(new_n390), .B2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(G20), .A2(G179), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT100), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT100), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n240), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n204), .A2(G190), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n398), .A3(new_n395), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G159), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n395), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n787), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(G20), .A3(G190), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n376), .B1(new_n793), .B2(new_n238), .C1(new_n527), .C2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n786), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n780), .B(KEYINPUT98), .Z(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n390), .A3(G200), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n390), .A3(new_n395), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n263), .A2(new_n798), .B1(new_n799), .B2(new_n354), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n797), .A2(G190), .A3(new_n395), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G58), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n796), .B(new_n803), .C1(new_n315), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n794), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G303), .A2(new_n810), .B1(new_n789), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n273), .C1(new_n812), .C2(new_n793), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G294), .B2(new_n784), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT33), .B(G317), .Z(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n799), .B1(new_n798), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G322), .B2(new_n802), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT101), .B(G326), .Z(new_n819));
  OAI211_X1 g0619(.A(new_n814), .B(new_n818), .C1(new_n808), .C2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n809), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n773), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n777), .B1(new_n778), .B2(new_n821), .C1(new_n689), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n400), .A2(new_n687), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n368), .A2(new_n687), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n391), .B2(new_n396), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(new_n400), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n713), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n698), .B(new_n829), .C1(new_n662), .C2(new_n668), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n761), .B1(new_n833), .B2(new_n754), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n754), .B2(new_n833), .ZN(new_n835));
  INV_X1    g0635(.A(new_n799), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n802), .B1(new_n836), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n258), .B2(new_n798), .C1(new_n808), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n376), .B1(new_n788), .B2(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n794), .A2(new_n315), .B1(new_n793), .B2(new_n263), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(new_n784), .C2(G58), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n793), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n848), .A2(G87), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n794), .A2(new_n238), .B1(new_n788), .B2(new_n815), .ZN(new_n850));
  NOR4_X1   g0650(.A1(new_n786), .A2(new_n376), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n549), .A2(new_n799), .B1(new_n798), .B2(new_n812), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G294), .B2(new_n802), .ZN(new_n853));
  INV_X1    g0653(.A(G303), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n851), .B(new_n853), .C1(new_n854), .C2(new_n808), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n774), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n774), .A2(new_n771), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n764), .B1(new_n354), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n772), .C2(new_n829), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n835), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT103), .Z(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n472), .A2(new_n477), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  OAI211_X1 g0665(.A(G116), .B(new_n221), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OR3_X1    g0668(.A1(new_n709), .A2(new_n354), .A3(new_n425), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n315), .A2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n203), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n440), .A2(new_n681), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n460), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n440), .A2(new_n441), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n873), .A3(new_n455), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n875), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n674), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n457), .A2(KEYINPUT104), .A3(new_n458), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n672), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n881), .B(new_n886), .C1(KEYINPUT38), .C2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n884), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n344), .A2(new_n686), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n672), .A2(new_n681), .ZN(new_n898));
  INV_X1    g0698(.A(new_n826), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n832), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n324), .A2(new_n687), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n343), .A2(new_n347), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n341), .A2(new_n340), .A3(G169), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n335), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n324), .B(new_n687), .C1(new_n905), .C2(new_n348), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n875), .A2(new_n880), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n881), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n898), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n897), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n461), .A2(new_n715), .A3(new_n719), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n676), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(G330), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n721), .B1(new_n569), .B2(new_n570), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n738), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n923), .A2(new_n830), .A3(new_n908), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n881), .B1(KEYINPUT38), .B2(new_n891), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT40), .B1(new_n912), .B2(new_n881), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n403), .A2(new_n460), .A3(new_n923), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n919), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n918), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n203), .B2(new_n758), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n918), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n872), .B1(new_n935), .B2(new_n936), .ZN(G367));
  NAND2_X1  g0737(.A1(new_n699), .A2(new_n487), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n521), .A2(new_n938), .A3(new_n525), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n663), .A2(new_n487), .A3(new_n699), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n697), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n521), .B1(new_n939), .B2(new_n613), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n942), .A2(KEYINPUT42), .B1(new_n698), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n563), .A2(new_n687), .ZN(new_n948));
  MUX2_X1   g0748(.A(new_n559), .B(new_n658), .S(new_n948), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT106), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n952), .A2(KEYINPUT107), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT107), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(KEYINPUT108), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n952), .A2(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT108), .B1(new_n955), .B2(new_n956), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n941), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n695), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n959), .A2(new_n963), .A3(new_n960), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n705), .B(KEYINPUT41), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n701), .A2(new_n941), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT45), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n701), .C2(new_n941), .ZN(new_n971));
  AND2_X1   g0771(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n972));
  NOR2_X1   g0772(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n973));
  OR4_X1    g0773(.A1(new_n701), .A2(new_n941), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n691), .A3(new_n694), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n695), .A3(new_n971), .A4(new_n974), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n696), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n619), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n694), .B2(new_n979), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n691), .B(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n720), .A2(new_n754), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n967), .B1(new_n985), .B2(new_n756), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n965), .A2(new_n966), .B1(new_n760), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n766), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n775), .B1(new_n207), .B2(new_n352), .C1(new_n988), .C2(new_n232), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n764), .B1(new_n989), .B2(KEYINPUT110), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT110), .B2(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT46), .B1(new_n810), .B2(G116), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT111), .Z(new_n993));
  INV_X1    g0793(.A(G294), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n785), .A2(new_n238), .B1(new_n994), .B2(new_n798), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n810), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT112), .B(G317), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n789), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n848), .A2(G97), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n998), .A3(new_n273), .A4(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n812), .A2(new_n799), .B1(new_n801), .B2(new_n854), .ZN(new_n1001));
  NOR4_X1   g0801(.A1(new_n993), .A2(new_n995), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n815), .B2(new_n808), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n808), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(G143), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G58), .A2(new_n810), .B1(new_n789), .B2(G137), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT113), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n793), .A2(new_n354), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n273), .ZN(new_n1009));
  OAI211_X1 g0809(.A(KEYINPUT113), .B(new_n376), .C1(new_n793), .C2(new_n354), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n836), .A2(G50), .B1(new_n784), .B2(G68), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n798), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G150), .A2(new_n802), .B1(new_n1013), .B2(G159), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1005), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1003), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n991), .B1(new_n1017), .B2(new_n774), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n822), .B2(new_n949), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n987), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT114), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  OR2_X1    g0823(.A1(new_n694), .A2(new_n822), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n766), .B1(new_n229), .B2(new_n290), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n768), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n707), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n256), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n707), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1027), .A2(new_n1031), .B1(new_n238), .B2(new_n704), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n775), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n761), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1004), .A2(G159), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n789), .A2(G150), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n810), .A2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n999), .A4(new_n376), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G68), .B2(new_n836), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n802), .A2(G50), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n785), .A2(new_n352), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n256), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n1013), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n819), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n376), .B1(new_n1045), .B2(new_n789), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n854), .A2(new_n799), .B1(new_n798), .B2(new_n815), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n802), .B2(new_n997), .ZN(new_n1048));
  INV_X1    g0848(.A(G322), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n808), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n784), .A2(G283), .B1(G294), .B2(new_n810), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1046), .B1(new_n549), .B2(new_n793), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1044), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1034), .B1(new_n1059), .B2(new_n774), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n982), .A2(new_n760), .B1(new_n1024), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n756), .A2(new_n982), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n983), .A2(new_n705), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(G393));
  NAND3_X1  g0864(.A1(new_n976), .A2(KEYINPUT115), .A3(new_n977), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n977), .A2(KEYINPUT115), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n983), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n985), .A2(new_n1067), .A3(new_n705), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT117), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n759), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n988), .A2(new_n244), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n775), .B1(new_n240), .B2(new_n207), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n761), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT116), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n1004), .A2(G317), .B1(G311), .B2(new_n802), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G283), .A2(new_n810), .B1(new_n789), .B2(G322), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n376), .B1(new_n848), .B2(G107), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n854), .C2(new_n798), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n785), .A2(new_n549), .B1(new_n994), .B2(new_n799), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1004), .A2(G150), .B1(G159), .B2(new_n802), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n849), .A2(new_n273), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G68), .A2(new_n810), .B1(new_n789), .B2(G143), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n256), .C2(new_n799), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n785), .A2(new_n354), .B1(new_n315), .B2(new_n798), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1075), .B1(new_n1090), .B2(new_n774), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n962), .A2(new_n773), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1069), .B1(new_n1071), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1093), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1070), .A2(KEYINPUT117), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1068), .B1(new_n1094), .B2(new_n1096), .ZN(G390));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n376), .B1(new_n793), .B2(new_n315), .C1(new_n1098), .C2(new_n788), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n810), .A2(G150), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G137), .C2(new_n1013), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1004), .A2(G128), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n802), .A2(G132), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n836), .A2(new_n1105), .B1(new_n784), .B2(G159), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n785), .A2(new_n354), .B1(new_n549), .B2(new_n801), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT121), .Z(new_n1109));
  AOI22_X1  g0909(.A1(G87), .A2(new_n810), .B1(new_n789), .B2(G294), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n376), .B1(new_n848), .B2(G68), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n240), .C2(new_n799), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G107), .B2(new_n1013), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n812), .B2(new_n808), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1107), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n778), .B1(new_n1115), .B2(KEYINPUT122), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n764), .B(new_n1119), .C1(new_n256), .C2(new_n858), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n895), .B2(new_n771), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n892), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n886), .B1(new_n912), .B2(new_n881), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT105), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n896), .B1(new_n900), .B2(new_n908), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n828), .A2(new_n400), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n686), .B(new_n1129), .C1(new_n718), .C2(new_n662), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n907), .B1(new_n1131), .B2(new_n826), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n896), .A3(new_n925), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n753), .A2(G330), .A3(new_n829), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(new_n908), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n829), .A2(new_n907), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(G330), .C1(new_n920), .C2(new_n922), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1122), .B1(new_n1140), .B2(new_n760), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(KEYINPUT120), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1138), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT120), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n923), .A2(new_n919), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n461), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n916), .A2(new_n676), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1134), .A2(new_n908), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1138), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n900), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT118), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT118), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1144), .B1(new_n1134), .B2(new_n908), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n900), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1150), .A2(new_n829), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n908), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1135), .A2(new_n1162), .A3(new_n899), .A4(new_n1130), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1152), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1142), .A2(new_n1149), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n705), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT118), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1158), .A2(new_n900), .A3(new_n1157), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1152), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1170), .A2(new_n1146), .A3(new_n1145), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT119), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT119), .B1(new_n1164), .B2(new_n1140), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1141), .B1(new_n1167), .B2(new_n1176), .ZN(G378));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n266), .A2(new_n681), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n312), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n312), .A2(new_n1180), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n926), .A2(KEYINPUT40), .B1(new_n924), .B2(new_n928), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n919), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n930), .A2(G330), .A3(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n915), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n897), .A2(new_n1190), .A3(new_n1191), .A4(new_n914), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1188), .A2(new_n771), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n774), .A2(G50), .A3(new_n771), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n376), .A2(G41), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G50), .B(new_n1198), .C1(new_n548), .C2(new_n289), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1004), .A2(G116), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G283), .A2(new_n789), .B1(new_n848), .B2(G58), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1037), .A3(new_n1198), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G68), .B2(new_n784), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n802), .A2(G107), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G97), .A2(new_n1013), .B1(new_n836), .B2(new_n366), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1200), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1199), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n843), .A2(new_n798), .B1(new_n799), .B2(new_n838), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G128), .B2(new_n802), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n784), .A2(G150), .B1(new_n810), .B2(new_n1105), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n1098), .C2(new_n808), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n848), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1208), .B1(new_n1207), .B2(new_n1206), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n764), .B(new_n1197), .C1(new_n1218), .C2(new_n774), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1195), .A2(new_n760), .B1(new_n1196), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1221), .B2(new_n1195), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1164), .A2(new_n1140), .A3(KEYINPUT119), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1152), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1195), .A2(KEYINPUT57), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n705), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1220), .B1(new_n1222), .B2(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n1170), .A2(new_n760), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n764), .B1(new_n263), .B2(new_n858), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n794), .A2(new_n240), .B1(new_n788), .B2(new_n854), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1041), .A2(new_n376), .A3(new_n1008), .A4(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n238), .A2(new_n799), .B1(new_n798), .B2(new_n549), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G283), .B2(new_n802), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n994), .C2(new_n808), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n808), .A2(new_n843), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G128), .A2(new_n789), .B1(new_n810), .B2(G159), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1238), .B(new_n376), .C1(new_n424), .C2(new_n793), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G150), .B2(new_n836), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1013), .A2(new_n1105), .B1(new_n784), .B2(G50), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n838), .C2(new_n801), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1236), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1231), .B1(new_n1243), .B2(new_n774), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n907), .B2(new_n772), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1229), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1164), .A2(new_n967), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1170), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1152), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(G381));
  NOR2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n862), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G390), .B1(KEYINPUT124), .B2(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1250), .A3(new_n1255), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G387), .A2(G378), .A3(G375), .A4(new_n1256), .ZN(G407));
  INV_X1    g1057(.A(new_n1141), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1164), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n706), .B1(new_n1259), .B2(new_n1142), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n683), .A2(new_n684), .A3(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G375), .C2(new_n1265), .ZN(G409));
  NAND2_X1  g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1268), .B2(new_n1252), .ZN(new_n1269));
  OR2_X1    g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1267), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G390), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1021), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(G390), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1020), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1020), .B(new_n1274), .C1(G390), .C2(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1220), .C1(new_n1222), .C2(new_n1227), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1195), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1225), .A2(new_n967), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1220), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1262), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1249), .A2(KEYINPUT60), .ZN(new_n1287));
  OR3_X1    g1087(.A1(new_n1170), .A2(KEYINPUT60), .A3(new_n1171), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1164), .A2(new_n706), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(new_n862), .A3(new_n1229), .A4(new_n1245), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1290), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1294));
  OAI21_X1  g1094(.A(G384), .B1(new_n1294), .B2(new_n1246), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1286), .A2(new_n1263), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1264), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(KEYINPUT125), .A3(new_n1296), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  XOR2_X1   g1102(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1303));
  NAND2_X1  g1103(.A1(new_n1286), .A2(new_n1263), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1264), .A2(G2897), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1296), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1292), .A2(new_n1295), .A3(new_n1305), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1303), .B1(new_n1304), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1280), .B1(new_n1302), .B2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(KEYINPUT61), .B(new_n1280), .C1(new_n1304), .C2(new_n1309), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1299), .A2(new_n1315), .A3(new_n1301), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1262), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1281), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1281), .A3(new_n1296), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XOR2_X1   g1124(.A(new_n1324), .B(new_n1280), .Z(G402));
endmodule


