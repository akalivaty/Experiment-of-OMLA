//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(G244), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(G77), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT16), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT7), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n248), .B1(new_n253), .B2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n248), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT74), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n249), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n258));
  AOI21_X1  g0058(.A(G33), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n203), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G58), .A2(G68), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n214), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G159), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(G20), .A3(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n247), .B1(new_n261), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n217), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n275), .A2(new_n276), .A3(new_n251), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n248), .B(new_n208), .C1(new_n277), .C2(new_n250), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G68), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n257), .A2(G33), .A3(new_n258), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n281));
  AOI21_X1  g0081(.A(G20), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n248), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n267), .B2(new_n270), .ZN(new_n285));
  AOI211_X1 g0085(.A(KEYINPUT76), .B(new_n269), .C1(new_n266), .C2(G20), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n279), .A2(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n272), .B(new_n274), .C1(new_n287), .C2(new_n247), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G13), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n296), .A2(new_n208), .A3(G1), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n274), .ZN(new_n298));
  INV_X1    g0098(.A(new_n292), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G223), .A2(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n280), .A3(new_n281), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G274), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n312), .B1(G232), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(G179), .ZN(new_n317));
  INV_X1    g0117(.A(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(G232), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n217), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G41), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n305), .B2(new_n306), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT77), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT77), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n309), .A2(new_n326), .A3(new_n315), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n317), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n301), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT18), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n288), .A2(new_n300), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n316), .A2(G190), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(KEYINPUT17), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G200), .B1(new_n325), .B2(new_n327), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n288), .B(new_n300), .C1(new_n340), .C2(new_n336), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n301), .A2(new_n330), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n332), .A2(new_n339), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n249), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n281), .A2(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n348), .A2(new_n303), .A3(G1698), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n281), .A2(new_n347), .A3(G232), .A4(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n308), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n310), .B1(new_n321), .B2(new_n322), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n314), .A2(G238), .B1(new_n355), .B2(new_n313), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n353), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g0159(.A(G169), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n360), .A2(KEYINPUT14), .B1(new_n361), .B2(G179), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(G169), .C1(new_n358), .C2(new_n359), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n356), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n329), .B1(new_n368), .B2(new_n357), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT73), .B1(new_n369), .B2(new_n363), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n362), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n298), .A2(G68), .A3(new_n293), .ZN(new_n372));
  XOR2_X1   g0172(.A(new_n372), .B(KEYINPUT72), .Z(new_n373));
  NOR2_X1   g0173(.A1(G20), .A2(G33), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n251), .A2(G20), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G77), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(new_n274), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n297), .A2(new_n203), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(KEYINPUT11), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n373), .A2(new_n381), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n385), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n368), .A2(new_n357), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n361), .A2(G190), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n293), .A2(G50), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n293), .A2(KEYINPUT68), .A3(G50), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n298), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n297), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(G50), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n274), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n292), .A2(new_n376), .B1(G150), .B2(new_n374), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n204), .A2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n312), .B1(G226), .B2(new_n314), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n281), .A2(new_n347), .A3(G222), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT66), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n348), .A2(G77), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n281), .A2(new_n347), .A3(G223), .A4(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT67), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n323), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT67), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n407), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n405), .B1(new_n423), .B2(G169), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT69), .ZN(new_n425));
  INV_X1    g0225(.A(new_n422), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n308), .B1(new_n421), .B2(KEYINPUT67), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n406), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n425), .B1(new_n428), .B2(G179), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(KEYINPUT69), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G232), .A2(G1698), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n408), .A2(G238), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n253), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n308), .C1(G107), .C2(new_n253), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n312), .B1(new_n220), .B2(new_n314), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G200), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n438), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n298), .A2(G77), .A3(new_n293), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT70), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n292), .A2(new_n374), .B1(G20), .B2(G77), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n377), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n274), .B1(new_n378), .B2(new_n297), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n438), .A2(new_n329), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n450), .C1(G179), .C2(new_n438), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n432), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT10), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n404), .A2(KEYINPUT9), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT9), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n399), .B2(new_n403), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(G200), .B2(new_n428), .ZN(new_n459));
  OAI211_X1 g0259(.A(G190), .B(new_n406), .C1(new_n426), .C2(new_n427), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n454), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n458), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n460), .C1(new_n423), .C2(new_n334), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT10), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n453), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(KEYINPUT71), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(KEYINPUT71), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n346), .B(new_n392), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n297), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(KEYINPUT25), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(KEYINPUT25), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n298), .B1(G1), .B2(new_n251), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n469), .ZN(new_n474));
  INV_X1    g0274(.A(G87), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n348), .A2(KEYINPUT22), .A3(G20), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n280), .A2(new_n208), .A3(G87), .A4(new_n281), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n478), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT84), .B1(new_n478), .B2(KEYINPUT22), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT81), .A2(G116), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT81), .A2(G116), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n251), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n208), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n469), .A2(G20), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT23), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT85), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n400), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n478), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n476), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n494), .B1(new_n499), .B2(new_n489), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n481), .A2(KEYINPUT85), .A3(new_n490), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(KEYINPUT24), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n474), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n280), .A2(new_n281), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G1698), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G250), .B2(G1698), .ZN(new_n507));
  INV_X1    g0307(.A(G294), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n504), .A2(new_n507), .B1(new_n251), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT79), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT78), .ZN(new_n511));
  INV_X1    g0311(.A(G41), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  INV_X1    g0313(.A(G45), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G1), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT78), .B1(new_n516), .B2(G41), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(G41), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n513), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n323), .A2(G274), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n511), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n516), .B2(G41), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n207), .A2(G45), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n518), .B2(new_n511), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n523), .A2(new_n525), .A3(new_n355), .A4(KEYINPUT79), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n509), .A2(new_n308), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n519), .A2(G264), .A3(new_n323), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(KEYINPUT86), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n519), .A2(new_n532), .A3(G264), .A4(new_n323), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n530), .B1(new_n430), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n503), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n474), .ZN(new_n539));
  AOI21_X1  g0339(.A(G200), .B1(new_n527), .B2(new_n534), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n509), .A2(new_n308), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n521), .A2(new_n526), .ZN(new_n542));
  AND4_X1   g0342(.A1(new_n440), .A2(new_n541), .A3(new_n542), .A4(new_n528), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n493), .B2(new_n502), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n473), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n482), .A2(new_n483), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(G116), .B1(new_n297), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n208), .C1(G33), .C2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n274), .B(new_n553), .C1(new_n548), .C2(new_n208), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n505), .A2(new_n408), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G264), .B2(new_n408), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n504), .A2(new_n559), .B1(new_n560), .B2(new_n253), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n308), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n519), .A2(G270), .A3(new_n323), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n542), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n557), .B1(G200), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n440), .B2(new_n564), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(new_n564), .A3(G169), .ZN(new_n567));
  NOR2_X1   g0367(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n568), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n557), .A2(new_n564), .A3(G169), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n564), .A2(new_n430), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n557), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n566), .A2(new_n569), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n445), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n398), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n473), .A2(new_n475), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n376), .A2(new_n578), .A3(G97), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n475), .B1(new_n351), .B2(new_n208), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(new_n581), .B2(new_n578), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n280), .A2(new_n208), .A3(G68), .A4(new_n281), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n400), .B1(new_n584), .B2(KEYINPUT82), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  AOI211_X1 g0387(.A(new_n576), .B(new_n577), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G238), .A2(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(G244), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(G1698), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n280), .A3(new_n281), .ZN(new_n592));
  INV_X1    g0392(.A(new_n484), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n323), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n524), .A2(G250), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n323), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n520), .B2(new_n524), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n594), .A2(new_n597), .A3(new_n440), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n355), .A2(new_n515), .B1(new_n595), .B2(new_n323), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n275), .A2(new_n276), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n250), .B1(new_n600), .B2(G33), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n484), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n599), .B1(new_n602), .B2(new_n323), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n598), .B1(G200), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n584), .A2(KEYINPUT82), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n274), .A3(new_n587), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n547), .A2(new_n575), .ZN(new_n607));
  INV_X1    g0407(.A(new_n576), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n430), .B(new_n599), .C1(new_n602), .C2(new_n323), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n329), .B1(new_n594), .B2(new_n597), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n588), .A2(new_n604), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n469), .B1(new_n254), .B2(new_n260), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n374), .A2(G77), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(new_n552), .A3(G107), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n208), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n274), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n398), .A2(G97), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n547), .B2(G97), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n590), .A2(G1698), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n504), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n281), .A2(new_n347), .A3(G250), .A4(G1698), .ZN(new_n630));
  AND2_X1   g0430(.A1(KEYINPUT4), .A2(G244), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n281), .A2(new_n347), .A3(new_n631), .A4(new_n408), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n630), .A2(new_n632), .A3(new_n551), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n308), .B1(new_n521), .B2(new_n526), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n519), .A2(G257), .A3(new_n323), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT80), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT80), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n519), .A2(new_n638), .A3(G257), .A4(new_n323), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(G200), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT4), .B1(new_n601), .B2(new_n627), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n630), .A2(new_n632), .A3(new_n551), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n308), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n440), .A2(new_n644), .A3(new_n640), .A4(new_n542), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n625), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n640), .A3(new_n430), .A4(new_n542), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n644), .A2(new_n640), .A3(new_n542), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n624), .B(new_n647), .C1(new_n648), .C2(G169), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n613), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n574), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n468), .A2(new_n546), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n544), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n500), .A2(KEYINPUT24), .A3(new_n501), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n274), .B1(new_n500), .B2(KEYINPUT24), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n624), .A2(new_n647), .ZN(new_n659));
  AOI21_X1  g0459(.A(G169), .B1(new_n635), .B2(new_n640), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n644), .A2(new_n640), .A3(new_n542), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n334), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n635), .A2(new_n440), .A3(new_n640), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n624), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n657), .A2(new_n658), .A3(new_n666), .A4(new_n613), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT87), .B1(new_n650), .B2(new_n545), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n503), .B2(new_n537), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n667), .A2(new_n668), .A3(new_n670), .A4(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n588), .A2(new_n604), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n609), .A2(new_n612), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n678), .B2(new_n649), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n613), .A2(new_n661), .A3(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n672), .A2(new_n674), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n468), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n386), .A2(new_n451), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n341), .B(KEYINPUT17), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(new_n391), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n301), .A2(new_n330), .A3(new_n344), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n344), .B1(new_n301), .B2(new_n330), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT89), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n464), .B2(new_n461), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n463), .A2(KEYINPUT10), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n459), .A2(new_n454), .A3(new_n460), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(KEYINPUT89), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n432), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n685), .A2(new_n699), .ZN(G369));
  INV_X1    g0500(.A(new_n669), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(G213), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT90), .Z(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(new_n557), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n574), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n546), .ZN(new_n715));
  INV_X1    g0515(.A(new_n709), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n503), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n538), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n715), .A2(new_n717), .B1(new_n718), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n669), .A2(new_n709), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n546), .A2(new_n721), .B1(new_n538), .B2(new_n716), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(G399));
  NAND3_X1  g0523(.A1(new_n211), .A2(KEYINPUT91), .A3(new_n512), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT91), .B1(new_n211), .B2(new_n512), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n580), .A2(new_n475), .A3(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n727), .A2(new_n207), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n216), .B2(new_n727), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n670), .A2(new_n657), .A3(new_n666), .A4(new_n613), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n709), .B1(new_n683), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n682), .B1(new_n671), .B2(KEYINPUT88), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n709), .B1(new_n736), .B2(new_n674), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n737), .B2(KEYINPUT29), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n546), .A2(new_n651), .A3(new_n716), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n594), .A2(new_n597), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(new_n534), .A3(new_n541), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n572), .A2(new_n741), .A3(new_n648), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n572), .A2(new_n741), .A3(new_n648), .A4(KEYINPUT30), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n740), .A2(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n662), .A2(new_n535), .A3(new_n746), .A4(new_n564), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n748), .B2(new_n709), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n738), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n732), .B1(new_n754), .B2(new_n207), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT92), .ZN(G364));
  INV_X1    g0556(.A(new_n727), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n296), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n207), .B1(new_n758), .B2(G45), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n211), .A2(new_n253), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n211), .ZN(new_n764));
  INV_X1    g0564(.A(new_n211), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n601), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n514), .B2(new_n216), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n242), .A2(new_n514), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n217), .B1(G20), .B2(new_n329), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n761), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n208), .A2(new_n430), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n440), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n348), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n208), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n782), .B(new_n786), .C1(G329), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n778), .A2(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n440), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G326), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(G190), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(G303), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n208), .B1(new_n779), .B2(new_n430), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(new_n440), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G294), .A2(new_n800), .B1(new_n802), .B2(G283), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n790), .A2(new_n793), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n788), .A2(new_n268), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  INV_X1    g0606(.A(new_n780), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n348), .B1(new_n807), .B2(G58), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(new_n378), .C2(new_n784), .ZN(new_n809));
  INV_X1    g0609(.A(new_n792), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n810), .A2(new_n201), .B1(new_n801), .B2(new_n469), .ZN(new_n811));
  INV_X1    g0611(.A(new_n794), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n203), .B1(new_n796), .B2(new_n475), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n809), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n799), .B(KEYINPUT93), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n552), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n804), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n777), .B1(new_n818), .B2(new_n774), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n773), .B(KEYINPUT94), .Z(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n712), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n713), .A2(new_n760), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n712), .A2(G330), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n452), .A2(new_n709), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n684), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n451), .A2(new_n709), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n709), .A2(new_n448), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n449), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n451), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n829), .B1(new_n737), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n753), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT99), .Z(new_n837));
  AOI21_X1  g0637(.A(new_n761), .B1(new_n835), .B2(new_n753), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n774), .A2(new_n771), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n760), .B1(new_n378), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G294), .A2(new_n807), .B1(new_n789), .B2(G311), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n348), .C1(new_n549), .C2(new_n784), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n810), .A2(new_n560), .B1(new_n796), .B2(new_n469), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n812), .A2(new_n845), .B1(new_n801), .B2(new_n475), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n817), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n784), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n807), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n810), .B2(new_n850), .C1(new_n851), .C2(new_n812), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  INV_X1    g0653(.A(KEYINPUT98), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n801), .A2(new_n203), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n797), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT97), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n504), .B1(G132), .B2(new_n789), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n202), .C2(new_n799), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n854), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n774), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n841), .B1(new_n862), .B2(new_n863), .C1(new_n772), .C2(new_n834), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n839), .A2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n758), .A2(new_n207), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n274), .B1(new_n287), .B2(new_n247), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n285), .A2(new_n286), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT7), .B1(new_n601), .B2(G20), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G68), .A3(new_n278), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n300), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n333), .A2(new_n338), .B1(new_n874), .B2(new_n706), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n330), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n301), .A2(new_n706), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n331), .A2(new_n878), .A3(new_n868), .A4(new_n341), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n706), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n687), .B2(new_n691), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n867), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n341), .ZN(new_n885));
  INV_X1    g0685(.A(new_n876), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n879), .ZN(new_n888));
  INV_X1    g0688(.A(new_n882), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n346), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n709), .A2(new_n385), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n369), .A2(new_n363), .B1(new_n388), .B2(new_n430), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n364), .A2(new_n365), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n369), .A2(KEYINPUT73), .A3(new_n363), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n391), .B(new_n893), .C1(new_n897), .C2(new_n387), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n385), .B(new_n709), .C1(new_n371), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT100), .B1(new_n829), .B2(new_n830), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT100), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n903), .B(new_n831), .C1(new_n684), .C2(new_n828), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n892), .B(new_n901), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n691), .A2(new_n706), .ZN(new_n906));
  INV_X1    g0706(.A(new_n878), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n346), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n331), .A2(new_n878), .A3(new_n341), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n879), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT102), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT39), .B1(new_n892), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n916), .A2(KEYINPUT102), .A3(new_n917), .A4(new_n891), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n386), .A2(new_n709), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n906), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n468), .B(new_n735), .C1(KEYINPUT29), .C2(new_n737), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n699), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(G330), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n468), .A2(new_n752), .ZN(new_n927));
  INV_X1    g0727(.A(new_n834), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n898), .B2(new_n900), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n930));
  INV_X1    g0730(.A(new_n913), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n908), .B2(new_n911), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n929), .B(new_n752), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT40), .B1(new_n884), .B2(new_n891), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n901), .A2(new_n834), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n739), .B2(new_n751), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n933), .A2(KEYINPUT40), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n926), .B1(new_n927), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n927), .B2(new_n938), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n866), .B1(new_n925), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n925), .B2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(new_n619), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n218), .A4(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n216), .A2(G77), .A3(new_n264), .A4(new_n265), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n203), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n296), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n766), .A2(new_n238), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n776), .B1(new_n765), .B2(new_n575), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n760), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n613), .B1(new_n716), .B2(new_n588), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n716), .A2(new_n588), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n677), .ZN(new_n957));
  NAND2_X1  g0757(.A1(KEYINPUT46), .A2(G116), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n812), .A2(new_n508), .B1(new_n796), .B2(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n810), .A2(new_n785), .B1(new_n801), .B2(new_n552), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n549), .B2(new_n796), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n780), .A2(new_n560), .B1(new_n784), .B2(new_n845), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G317), .B2(new_n789), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n601), .B1(G107), .B2(new_n800), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n961), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n796), .A2(new_n202), .B1(new_n788), .B2(new_n850), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT110), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n815), .A2(G68), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n253), .B1(new_n780), .B2(new_n851), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G50), .B2(new_n848), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n792), .A2(G143), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n794), .A2(G159), .B1(new_n802), .B2(G77), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n967), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT111), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  OAI221_X1 g0778(.A(new_n954), .B1(new_n820), .B2(new_n957), .C1(new_n978), .C2(new_n863), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT112), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n546), .A2(new_n721), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n666), .B1(new_n625), .B2(new_n716), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n661), .A2(new_n709), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT103), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n649), .B1(new_n718), .B2(new_n982), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n987), .A2(KEYINPUT42), .B1(new_n716), .B2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(new_n991), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n720), .A2(new_n985), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n759), .B(KEYINPUT107), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n722), .A2(new_n984), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n720), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(KEYINPUT106), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n722), .A2(new_n984), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT105), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1003), .B2(KEYINPUT105), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1002), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n754), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n981), .B1(new_n719), .B2(new_n721), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n714), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n754), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n727), .B(KEYINPUT41), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n998), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n996), .A2(KEYINPUT108), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT108), .B1(new_n996), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n980), .B1(new_n1020), .B2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n1014), .A2(new_n997), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G303), .A2(new_n848), .B1(new_n807), .B2(G317), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n810), .B2(new_n781), .C1(new_n785), .C2(new_n812), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G283), .A2(new_n800), .B1(new_n797), .B2(G294), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT49), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n601), .B1(G326), .B2(new_n789), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n549), .B2(new_n801), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n815), .A2(new_n575), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n810), .A2(new_n268), .B1(new_n796), .B2(new_n378), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n292), .B2(new_n794), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n784), .A2(new_n203), .B1(new_n788), .B2(new_n851), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G50), .B2(new_n807), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n504), .B1(G97), .B2(new_n802), .ZN(new_n1040));
  AND4_X1   g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n774), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n729), .C1(G68), .C2(G77), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n299), .B2(G50), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n299), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n766), .C1(new_n235), .C2(new_n514), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n729), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(G107), .B2(new_n211), .C1(new_n1050), .C2(new_n762), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n760), .B1(new_n1051), .B2(new_n775), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1042), .B(new_n1052), .C1(new_n719), .C2(new_n820), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1015), .A2(new_n727), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1023), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(G393));
  AOI21_X1  g0856(.A(new_n757), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n985), .A2(new_n773), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n775), .B1(new_n552), .B2(new_n211), .C1(new_n767), .C2(new_n245), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n761), .A2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n810), .A2(new_n851), .B1(new_n268), .B2(new_n780), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT51), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n815), .A2(G77), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n797), .A2(G68), .B1(new_n802), .B2(G87), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n292), .A2(new_n848), .B1(new_n789), .B2(G143), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n794), .A2(G50), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n601), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n792), .A2(G317), .B1(new_n807), .B2(G311), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n812), .A2(new_n560), .B1(new_n801), .B2(new_n469), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n348), .B1(new_n788), .B2(new_n781), .C1(new_n508), .C2(new_n784), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n549), .A2(new_n799), .B1(new_n796), .B2(new_n845), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1067), .A2(new_n1071), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n774), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1011), .A2(new_n997), .B1(new_n1059), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1058), .A2(new_n1080), .ZN(G390));
  NOR2_X1   g0881(.A1(new_n753), .A2(new_n928), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n901), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n920), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n919), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n833), .A2(new_n451), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n831), .B1(new_n734), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n901), .B(KEYINPUT114), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n916), .A2(new_n891), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1086), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1084), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1094), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n829), .A2(KEYINPUT100), .A3(new_n830), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n828), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n736), .B2(new_n674), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n903), .B1(new_n1099), .B2(new_n831), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n920), .B1(new_n1101), .B2(new_n901), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1083), .B(new_n1096), .C1(new_n1102), .C2(new_n919), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n468), .A2(G330), .A3(new_n752), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n923), .A2(new_n699), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1082), .A2(new_n901), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1101), .B1(new_n1084), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1090), .B1(new_n753), .B2(new_n928), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1083), .A2(new_n1089), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1095), .A2(new_n1103), .A3(new_n1111), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n727), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1095), .A2(new_n1103), .A3(new_n997), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n840), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n761), .B1(new_n292), .B2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n784), .A2(new_n552), .B1(new_n788), .B2(new_n508), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n253), .B(new_n1119), .C1(G116), .C2(new_n807), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n855), .B1(G87), .B2(new_n797), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n794), .A2(G107), .B1(new_n792), .B2(G283), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1120), .A2(new_n1065), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n792), .A2(G128), .B1(new_n802), .B2(G50), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n850), .B2(new_n812), .C1(new_n816), .C2(new_n268), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n796), .A2(new_n851), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n848), .ZN(new_n1130));
  INV_X1    g0930(.A(G132), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n253), .B1(new_n780), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G125), .B2(new_n789), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1127), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1123), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1118), .B1(new_n1135), .B2(new_n774), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n919), .B2(new_n772), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1116), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1115), .A2(new_n1138), .ZN(G378));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n707), .A2(new_n404), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n432), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n698), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n432), .B(new_n1142), .C1(new_n694), .C2(new_n697), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n464), .A2(new_n461), .A3(new_n693), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT89), .B1(new_n695), .B2(new_n696), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1144), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1142), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n698), .A2(new_n1144), .A3(new_n1143), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n1140), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1147), .A2(new_n1153), .A3(KEYINPUT118), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n937), .B2(new_n926), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1147), .A2(new_n1153), .A3(KEYINPUT118), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n934), .A2(new_n936), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT40), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n936), .B2(new_n1092), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1156), .B(G330), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n905), .A2(new_n1155), .A3(new_n921), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n905), .A2(new_n921), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n997), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1147), .A2(new_n1153), .A3(new_n771), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n760), .B1(new_n201), .B2(new_n840), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n807), .B1(new_n848), .B2(G137), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n792), .A2(G125), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n1131), .C2(new_n812), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1129), .A2(new_n797), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n816), .A2(new_n851), .B1(new_n1172), .B2(KEYINPUT116), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(KEYINPUT116), .C2(new_n1172), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n802), .A2(G159), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G107), .A2(new_n807), .B1(new_n848), .B2(new_n575), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n845), .B2(new_n788), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n552), .A2(new_n812), .B1(new_n810), .B2(new_n728), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n202), .A2(new_n801), .B1(new_n796), .B2(new_n378), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n601), .A2(G41), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1187), .A2(new_n970), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1191));
  AND4_X1   g0991(.A1(new_n1180), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1167), .B(new_n1168), .C1(new_n863), .C2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT117), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1166), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1106), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1197), .C1(new_n1198), .C2(new_n1114), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1114), .A2(new_n1198), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1197), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT119), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1165), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n757), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1195), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G375));
  INV_X1    g1008(.A(new_n1018), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1112), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n998), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1090), .A2(new_n771), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n761), .B1(G68), .B2(new_n1117), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n796), .A2(new_n552), .B1(new_n788), .B2(new_n560), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT120), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n348), .B1(new_n780), .B2(new_n845), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G107), .B2(new_n848), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n794), .A2(new_n548), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n792), .A2(G294), .B1(new_n802), .B2(G77), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1035), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n815), .A2(G50), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1129), .A2(new_n794), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n780), .A2(new_n850), .B1(new_n784), .B2(new_n851), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(new_n504), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n792), .A2(G132), .B1(new_n802), .B2(G58), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n797), .A2(G159), .B1(new_n789), .B2(G128), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT121), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1216), .A2(new_n1221), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1214), .B1(new_n1230), .B2(new_n774), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1212), .B1(new_n1213), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1211), .A2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(G390), .ZN(new_n1234));
  INV_X1    g1034(.A(G384), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1236), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1237));
  INV_X1    g1037(.A(G387), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1207), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n708), .A2(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1207), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  INV_X1    g1044(.A(KEYINPUT61), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1166), .A2(new_n1193), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1114), .A2(new_n1198), .B1(new_n1164), .B2(new_n1162), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n1209), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G378), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1207), .B2(G378), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT125), .B1(new_n1250), .B2(new_n1242), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1242), .A2(G2897), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1210), .B1(new_n1111), .B2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT60), .A4(new_n1110), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n727), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1258), .B(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(G384), .A3(new_n1232), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1260), .B2(new_n1232), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1254), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1232), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1235), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(G384), .A3(new_n1232), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1253), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1195), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1197), .B1(new_n1114), .B2(new_n1198), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT119), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n727), .B1(new_n1247), .B2(KEYINPUT57), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G378), .B(new_n1269), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1249), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1241), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1251), .A2(new_n1268), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1251), .B2(new_n1277), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1245), .B(new_n1278), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1275), .A2(KEYINPUT122), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1241), .B1(new_n1275), .B2(KEYINPUT122), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1284), .A2(new_n1285), .A3(KEYINPUT62), .A4(new_n1280), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1251), .A2(new_n1277), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT62), .B1(new_n1288), .B2(new_n1280), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1278), .A2(new_n1245), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1282), .A3(new_n1279), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(G393), .B(new_n826), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1234), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n980), .B(G390), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1287), .A2(new_n1294), .A3(new_n1303), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1284), .A2(new_n1285), .A3(new_n1280), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1305), .A2(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1281), .A2(KEYINPUT63), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1268), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(G405));
  XNOR2_X1  g1112(.A(new_n1207), .B(G378), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(new_n1279), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(new_n1307), .ZN(G402));
endmodule


