//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(new_n206), .A2(G50), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  NAND4_X1  g0013(.A1(new_n213), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G77), .Z(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n218), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n214), .B(new_n221), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n245), .B(new_n251), .Z(G351));
  OAI21_X1  g0052(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT8), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n257), .A2(KEYINPUT68), .A3(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n216), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n215), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n265), .A3(new_n264), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(new_n272), .B2(G50), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n286), .B1(new_n222), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n265), .B1(G33), .B2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  OAI211_X1 g0094(.A(G1), .B(G13), .C1(new_n281), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n295), .A3(G274), .ZN(new_n296));
  INV_X1    g0096(.A(G226), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n290), .A2(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n291), .B(new_n296), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n301), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n277), .B2(new_n278), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n279), .A2(new_n308), .B1(new_n310), .B2(new_n303), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n256), .A2(new_n246), .B1(new_n216), .B2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n262), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n266), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  INV_X1    g0120(.A(new_n268), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n203), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n203), .B2(new_n271), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G238), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n296), .B1(new_n327), .B2(new_n299), .C1(new_n331), .C2(new_n295), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(G169), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n333), .B2(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n326), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT72), .B1(new_n333), .B2(new_n305), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n332), .B(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(G190), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n326), .B1(new_n333), .B2(G200), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n300), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n274), .C1(G179), .C2(new_n300), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n296), .B1(new_n299), .B2(new_n223), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n284), .A2(G232), .A3(new_n285), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n353), .B1(new_n209), .B2(new_n284), .C1(new_n287), .C2(new_n327), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT69), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n295), .B1(new_n354), .B2(new_n355), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G179), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT15), .B(G87), .Z(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n362), .A2(new_n262), .B1(new_n216), .B2(new_n222), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n259), .A2(new_n256), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n266), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n272), .A2(G77), .B1(new_n222), .B2(new_n321), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n358), .B2(G169), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n358), .B2(G190), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n358), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n311), .A2(new_n348), .A3(new_n351), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n282), .A2(new_n216), .A3(new_n283), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT7), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n282), .A2(new_n377), .A3(new_n216), .A4(new_n283), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(G68), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G159), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n380), .A2(G20), .A3(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n204), .A2(new_n205), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n383), .B2(G20), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI211_X1 g0187(.A(new_n386), .B(new_n381), .C1(new_n383), .C2(G20), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n376), .B2(new_n378), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n203), .B1(new_n375), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n388), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(new_n394), .A3(new_n266), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n257), .A2(G58), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT68), .ZN(new_n399));
  OR3_X1    g0199(.A1(new_n257), .A2(KEYINPUT68), .A3(G58), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(new_n271), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n321), .B1(new_n399), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n271), .A3(new_n400), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(KEYINPUT74), .C1(new_n260), .C2(new_n321), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n288), .A2(new_n285), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n297), .A2(G1698), .ZN(new_n409));
  AND2_X1   g0209(.A1(KEYINPUT3), .A2(G33), .ZN(new_n410));
  NOR2_X1   g0210(.A1(KEYINPUT3), .A2(G33), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G87), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n281), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n295), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI211_X1 g0218(.A(KEYINPUT75), .B(new_n295), .C1(new_n412), .C2(new_n415), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n295), .A2(G232), .A3(new_n292), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n296), .A2(new_n420), .A3(new_n336), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n296), .A2(new_n420), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n416), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT76), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  INV_X1    g0227(.A(new_n421), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G223), .A2(G1698), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n297), .B2(G1698), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n414), .B1(new_n430), .B2(new_n284), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT75), .B1(new_n431), .B2(new_n295), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n416), .A2(new_n417), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n435), .C1(G169), .C2(new_n424), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n407), .A2(new_n426), .A3(new_n427), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n407), .A2(new_n426), .A3(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT18), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n296), .A2(new_n420), .A3(new_n305), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n432), .A2(new_n433), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n371), .B1(new_n423), .B2(new_n416), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n395), .A2(new_n443), .A3(new_n406), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n395), .A2(new_n443), .A3(new_n406), .A4(new_n445), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n437), .B(new_n439), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n374), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n284), .A2(G264), .A3(G1698), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(new_n285), .C1(new_n410), .C2(new_n411), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n410), .A2(new_n411), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G303), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n290), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT5), .B(G41), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n290), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G274), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n290), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n466), .A2(G270), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n266), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n215), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(G116), .A3(new_n268), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n264), .A2(new_n265), .B1(G20), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n216), .C1(G33), .C2(new_n208), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT20), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  OAI221_X1 g0283(.A(new_n477), .B1(G116), .B2(new_n268), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n474), .A2(new_n484), .A3(KEYINPUT21), .A4(G169), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n473), .A3(new_n462), .A4(G179), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n349), .B1(new_n462), .B2(new_n473), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT21), .B1(new_n488), .B2(new_n484), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n484), .B1(new_n474), .B2(G200), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n305), .B2(new_n474), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n465), .A2(new_n295), .A3(G274), .A4(new_n464), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n471), .A2(new_n295), .ZN(new_n495));
  INV_X1    g0295(.A(G257), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(new_n285), .C1(new_n410), .C2(new_n411), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n499), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n284), .A2(G244), .A3(new_n285), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n502), .A3(new_n480), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n497), .B1(new_n504), .B2(new_n290), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G190), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n321), .A2(new_n208), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n475), .A2(new_n268), .A3(new_n476), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n208), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n376), .A2(G107), .A3(new_n378), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n255), .A2(G77), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT79), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n209), .A2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n210), .A2(new_n513), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(G20), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n510), .A2(new_n511), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n509), .B1(new_n522), .B2(new_n266), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  OAI21_X1  g0324(.A(G200), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(KEYINPUT81), .B(new_n497), .C1(new_n290), .C2(new_n504), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n506), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G238), .B(new_n285), .C1(new_n410), .C2(new_n411), .ZN(new_n528));
  OAI211_X1 g0328(.A(G244), .B(G1698), .C1(new_n410), .C2(new_n411), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n290), .ZN(new_n532));
  INV_X1    g0332(.A(G250), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n464), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n468), .A2(new_n464), .B1(new_n534), .B2(new_n295), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n361), .A2(new_n268), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n268), .A2(new_n476), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n413), .A3(new_n266), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n216), .B1(new_n330), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n413), .A2(new_n208), .A3(new_n209), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n216), .B(G68), .C1(new_n410), .C2(new_n411), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n541), .B1(new_n262), .B2(new_n208), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n538), .B(new_n540), .C1(new_n266), .C2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n532), .A2(new_n535), .A3(G190), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n537), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n547), .B2(new_n266), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n508), .A2(new_n362), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n532), .A2(new_n535), .A3(new_n336), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n534), .A2(new_n295), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n295), .A2(G274), .A3(new_n464), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n290), .B2(new_n531), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(G169), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n504), .A2(new_n290), .ZN(new_n561));
  INV_X1    g0361(.A(new_n497), .ZN(new_n562));
  AOI21_X1  g0362(.A(G169), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n523), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n505), .A2(new_n336), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n527), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(G1698), .C1(new_n410), .C2(new_n411), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(new_n285), .C1(new_n410), .C2(new_n411), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G294), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n290), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n466), .A2(G264), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(G179), .A3(new_n494), .A4(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n471), .A2(new_n290), .A3(new_n467), .ZN(new_n580));
  OAI21_X1  g0380(.A(G169), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n216), .B(G87), .C1(new_n410), .C2(new_n411), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT22), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT22), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n284), .A2(new_n585), .A3(new_n216), .A4(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n530), .A2(G20), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n216), .A2(G107), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n590), .A2(KEYINPUT23), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(KEYINPUT23), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n587), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n588), .B1(new_n587), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n266), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G13), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(G1), .ZN(new_n598));
  OR2_X1    g0398(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n599));
  NAND2_X1  g0399(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n590), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n598), .A2(new_n590), .ZN(new_n602));
  OAI221_X1 g0402(.A(new_n601), .B1(new_n602), .B2(new_n600), .C1(new_n508), .C2(new_n209), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n582), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n576), .A2(new_n494), .A3(new_n578), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n371), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n573), .A2(new_n574), .A3(new_n305), .A4(new_n494), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR4_X1   g0411(.A1(new_n493), .A2(new_n568), .A3(new_n607), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n456), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n613), .B(KEYINPUT84), .Z(G372));
  NOR2_X1   g0414(.A1(new_n563), .A2(new_n523), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(new_n566), .A3(new_n559), .A4(new_n550), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT85), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n560), .A3(new_n620), .A4(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n606), .A2(new_n490), .ZN(new_n624));
  INV_X1    g0424(.A(new_n505), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n505), .A2(new_n524), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G200), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n506), .A2(new_n523), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(new_n629), .B1(new_n615), .B2(new_n566), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n577), .B1(new_n573), .B2(new_n574), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n631), .A2(new_n632), .A3(new_n580), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n610), .B1(new_n633), .B2(G200), .ZN(new_n634));
  INV_X1    g0434(.A(new_n605), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n624), .A2(new_n630), .A3(new_n560), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(new_n637), .A3(new_n559), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n456), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n369), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n347), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n403), .A2(new_n405), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n377), .B1(new_n459), .B2(new_n216), .ZN(new_n643));
  INV_X1    g0443(.A(new_n378), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT73), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n392), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n475), .B1(new_n646), .B2(new_n388), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n642), .B1(new_n647), .B2(new_n387), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n448), .B1(new_n648), .B2(new_n443), .ZN(new_n649));
  INV_X1    g0449(.A(new_n452), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT78), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n641), .A2(new_n339), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n422), .A2(new_n425), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n407), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(new_n427), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n311), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n351), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n639), .A2(new_n659), .ZN(G369));
  NAND2_X1  g0460(.A1(new_n598), .A2(new_n216), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n636), .B(new_n606), .C1(new_n635), .C2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT88), .Z(new_n669));
  NOR2_X1   g0469(.A1(new_n490), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n607), .A2(new_n667), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n484), .A2(new_n666), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n493), .B2(KEYINPUT86), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(KEYINPUT86), .B2(new_n493), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n490), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT87), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n606), .A2(new_n667), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n669), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n677), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n219), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n543), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n213), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n693), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n474), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(G179), .A3(new_n505), .A4(new_n558), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n700), .A2(new_n632), .A3(new_n631), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n699), .A2(G179), .A3(new_n558), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n625), .A3(new_n608), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n666), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n612), .A2(new_n667), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n559), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n568), .A2(new_n611), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n624), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n666), .B1(new_n717), .B2(new_n623), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n616), .B(new_n617), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n666), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(KEYINPUT29), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n698), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n597), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n215), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OR3_X1    g0527(.A1(new_n692), .A2(KEYINPUT90), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT90), .B1(new_n692), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n684), .B2(G330), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n684), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT91), .Z(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n683), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n265), .B1(G20), .B2(new_n349), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n213), .A2(new_n463), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n691), .A2(new_n284), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(new_n743), .C1(new_n463), .C2(new_n251), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n691), .A2(new_n459), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(G355), .B1(new_n478), .B2(new_n691), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n741), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n739), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n216), .A2(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT32), .B1(new_n751), .B2(new_n380), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n216), .A2(new_n336), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n305), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n752), .B1(new_n756), .B2(new_n246), .C1(new_n203), .C2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n216), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n208), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n751), .A2(KEYINPUT32), .A3(new_n380), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n413), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n749), .A2(new_n305), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n209), .ZN(new_n767));
  OR4_X1    g0567(.A1(new_n762), .A2(new_n763), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n753), .A2(new_n750), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n753), .A2(G190), .A3(new_n371), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n284), .B1(new_n222), .B2(new_n769), .C1(new_n202), .C2(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n759), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n766), .A2(new_n773), .B1(new_n751), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT92), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n459), .B1(new_n769), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n770), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G322), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n761), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G294), .A2(new_n781), .B1(new_n755), .B2(G326), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  INV_X1    g0583(.A(new_n764), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n757), .A2(new_n783), .B1(new_n784), .B2(G303), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n776), .A2(new_n780), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n748), .B1(new_n772), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n747), .A2(new_n787), .A3(new_n730), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n738), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n734), .A2(new_n789), .ZN(G396));
  NOR3_X1   g0590(.A1(new_n360), .A2(new_n368), .A3(new_n666), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n367), .A2(new_n666), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n372), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n793), .B2(new_n369), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT96), .ZN(new_n795));
  INV_X1    g0595(.A(new_n718), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n638), .A2(new_n667), .A3(new_n794), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n638), .A2(KEYINPUT97), .A3(new_n794), .A4(new_n667), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n731), .B1(new_n803), .B2(new_n713), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n713), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n739), .A2(new_n735), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n731), .B1(G77), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n769), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n755), .A2(G303), .B1(new_n809), .B2(G116), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n773), .B2(new_n758), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT93), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n766), .A2(new_n413), .B1(new_n751), .B2(new_n777), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n459), .B1(new_n770), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n762), .B(new_n816), .C1(G107), .C2(new_n784), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n812), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n779), .A2(G143), .B1(new_n809), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n756), .B2(new_n820), .C1(new_n254), .C2(new_n758), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  OAI22_X1  g0622(.A1(new_n246), .A2(new_n764), .B1(new_n766), .B2(new_n203), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT95), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n284), .B1(new_n751), .B2(new_n826), .C1(new_n761), .C2(new_n202), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n824), .B2(new_n823), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n818), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n808), .B1(new_n830), .B2(new_n739), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n794), .B2(new_n736), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n805), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(new_n222), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n213), .A2(new_n834), .A3(new_n382), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n215), .B(G13), .C1(new_n835), .C2(new_n247), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n265), .A2(new_n216), .A3(new_n478), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n518), .A2(new_n520), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT35), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT36), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(new_n664), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n407), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g0646(.A1(new_n844), .A2(new_n438), .A3(new_n444), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n404), .B1(new_n260), .B2(new_n321), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n646), .B2(new_n384), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n394), .A2(new_n266), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(KEYINPUT99), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n654), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n845), .A3(new_n854), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n444), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n847), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n651), .A2(new_n652), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n439), .A2(new_n437), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n856), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n856), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT100), .B1(new_n455), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(KEYINPUT38), .B(new_n859), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n655), .A2(new_n846), .A3(new_n444), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n847), .B1(KEYINPUT37), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n450), .A2(new_n452), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n846), .B1(new_n656), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n867), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n347), .ZN(new_n874));
  INV_X1    g0674(.A(new_n338), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(new_n335), .C1(new_n336), .C2(new_n333), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n326), .B(new_n666), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n339), .B(new_n347), .C1(new_n325), .C2(new_n667), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n712), .A3(new_n794), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n873), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n880), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n859), .B1(new_n863), .B2(new_n865), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n867), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(new_n886), .A3(new_n866), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n885), .B2(new_n866), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n882), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(new_n456), .A3(new_n712), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G330), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n456), .B2(new_n712), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n439), .A2(new_n437), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n651), .B2(new_n652), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n860), .B1(new_n896), .B2(new_n856), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n455), .A2(KEYINPUT100), .A3(new_n864), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n899), .B2(new_n859), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n867), .B(new_n858), .C1(new_n897), .C2(new_n898), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT101), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n885), .A2(new_n886), .A3(new_n866), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT98), .ZN(new_n906));
  INV_X1    g0706(.A(new_n791), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n802), .B2(new_n907), .ZN(new_n908));
  AOI211_X1 g0708(.A(KEYINPUT98), .B(new_n791), .C1(new_n800), .C2(new_n801), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n879), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n905), .A2(new_n910), .B1(new_n656), .B2(new_n845), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n876), .A2(new_n326), .A3(new_n667), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n885), .B2(new_n866), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n913), .B2(new_n873), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n900), .B2(new_n901), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT102), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n911), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n456), .A2(new_n722), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n659), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n894), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n215), .B2(new_n725), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n894), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n843), .B1(new_n925), .B2(new_n926), .ZN(G367));
  OAI21_X1  g0727(.A(new_n630), .B1(new_n523), .B2(new_n667), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n619), .A2(new_n666), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n689), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n560), .B1(new_n548), .B2(new_n667), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n559), .A2(new_n548), .A3(new_n667), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT43), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n669), .A2(new_n670), .A3(new_n930), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n607), .A2(new_n527), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n666), .B1(new_n944), .B2(new_n567), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n941), .B2(KEYINPUT42), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n940), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT43), .B2(new_n937), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n943), .A2(new_n939), .A3(new_n938), .A4(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n932), .A2(new_n933), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n933), .B(new_n932), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n692), .B(KEYINPUT41), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n931), .B1(new_n674), .B2(new_n676), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT45), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n674), .A2(new_n676), .A3(new_n931), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n688), .ZN(new_n962));
  INV_X1    g0762(.A(new_n687), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n671), .B1(new_n963), .B2(new_n670), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(new_n685), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n723), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n960), .A3(new_n689), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n962), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n955), .B1(new_n969), .B2(new_n723), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n954), .B1(new_n970), .B2(new_n727), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n938), .A2(new_n737), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n743), .A2(new_n241), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n741), .B1(new_n691), .B2(new_n361), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n730), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n766), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G159), .A2(new_n757), .B1(new_n834), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n202), .B2(new_n764), .ZN(new_n978));
  INV_X1    g0778(.A(new_n751), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n779), .A2(G150), .B1(new_n979), .B2(G137), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n284), .C1(new_n246), .C2(new_n769), .ZN(new_n981));
  INV_X1    g0781(.A(G143), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n756), .A2(new_n982), .B1(new_n203), .B2(new_n761), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT106), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n779), .A2(G303), .B1(new_n979), .B2(G317), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n459), .C1(new_n773), .C2(new_n769), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n764), .A2(new_n478), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(KEYINPUT46), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(KEYINPUT46), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT105), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G107), .A2(new_n781), .B1(new_n755), .B2(G311), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n757), .A2(G294), .B1(new_n976), .B2(G97), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n989), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI211_X1 g0796(.A(new_n972), .B(new_n975), .C1(new_n996), .C2(new_n748), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n971), .A2(new_n997), .ZN(G387));
  NAND2_X1  g0798(.A1(new_n687), .A2(new_n737), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n463), .B1(new_n203), .B2(new_n313), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n259), .A2(G50), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT108), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n743), .B1(new_n238), .B2(new_n463), .C1(new_n1005), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n694), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n745), .A2(new_n1011), .B1(new_n209), .B2(new_n691), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n741), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n459), .B1(new_n979), .B2(G150), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n208), .B2(new_n766), .C1(new_n222), .C2(new_n764), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT109), .Z(new_n1016));
  AOI22_X1  g0816(.A1(new_n779), .A2(G50), .B1(new_n809), .B2(G68), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n362), .B2(new_n761), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G159), .B2(new_n755), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(new_n261), .C2(new_n758), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n284), .B1(new_n979), .B2(G326), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n761), .A2(new_n773), .B1(new_n764), .B2(new_n815), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n779), .A2(G317), .B1(new_n809), .B2(G303), .ZN(new_n1023));
  INV_X1    g0823(.A(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(new_n756), .B2(new_n1024), .C1(new_n777), .C2(new_n758), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1021), .B1(new_n478), .B2(new_n766), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n730), .B(new_n1013), .C1(new_n1032), .C2(new_n739), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n965), .A2(new_n727), .B1(new_n999), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n966), .A2(new_n692), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n965), .A2(new_n723), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(G393));
  INV_X1    g0837(.A(new_n968), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n689), .B1(new_n957), .B2(new_n960), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n931), .A2(new_n737), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n740), .B1(new_n208), .B2(new_n219), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n743), .B2(new_n245), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT110), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G150), .A2(new_n755), .B1(new_n779), .B2(G159), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n758), .A2(new_n246), .B1(new_n766), .B2(new_n413), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n284), .B1(new_n751), .B2(new_n982), .C1(new_n259), .C2(new_n769), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n761), .A2(new_n313), .B1(new_n764), .B2(new_n203), .ZN(new_n1049));
  OR3_X1    g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n284), .B(new_n767), .C1(G294), .C2(new_n809), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n764), .A2(new_n773), .B1(new_n751), .B2(new_n1024), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT111), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(KEYINPUT111), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G116), .A2(new_n781), .B1(new_n757), .B2(G303), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n755), .B1(new_n779), .B2(G311), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1046), .A2(new_n1050), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n730), .B(new_n1044), .C1(new_n1059), .C2(new_n739), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT112), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1040), .A2(new_n727), .B1(new_n1041), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n966), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n969), .A3(new_n692), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(G390));
  NAND3_X1  g0865(.A1(new_n712), .A2(G330), .A3(new_n794), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n879), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n793), .A2(new_n369), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n791), .B1(new_n721), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n873), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n912), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n873), .A2(new_n913), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n915), .B(KEYINPUT39), .C1(new_n900), .C2(new_n901), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n914), .A2(new_n915), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n910), .A2(new_n912), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1068), .B(new_n1073), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1068), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT97), .B1(new_n718), .B2(new_n794), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n801), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n907), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT98), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n802), .A2(new_n906), .A3(new_n907), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n912), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n918), .B(new_n916), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1073), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1081), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1080), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n456), .A2(new_n714), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n921), .A2(new_n1093), .A3(new_n659), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1068), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1067), .B1(new_n713), .B2(new_n795), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1081), .A2(new_n1070), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n693), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1088), .B1(new_n1095), .B2(new_n879), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n918), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1090), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1068), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1089), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1100), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT113), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1110), .B(new_n1100), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1101), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n730), .B1(new_n261), .B2(new_n806), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n459), .B1(new_n979), .B2(G125), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n246), .B2(new_n766), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT115), .Z(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1117));
  NOR3_X1   g0917(.A1(new_n1117), .A2(new_n764), .A3(new_n254), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n764), .B2(new_n254), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n826), .B2(new_n770), .C1(new_n756), .C2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1116), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n781), .A2(G159), .B1(new_n809), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n820), .B2(new_n758), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT114), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n756), .A2(new_n773), .B1(new_n313), .B2(new_n761), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n459), .B1(new_n751), .B2(new_n815), .C1(new_n770), .C2(new_n478), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n766), .A2(new_n203), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1128), .A2(new_n765), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n757), .A2(G107), .B1(new_n809), .B2(G97), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT117), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1122), .A2(new_n1127), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1113), .B1(new_n748), .B2(new_n1134), .C1(new_n1103), .C2(new_n736), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1107), .B2(new_n726), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1112), .A2(new_n1137), .ZN(G378));
  OAI21_X1  g0938(.A(KEYINPUT120), .B1(new_n911), .B2(new_n919), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n275), .A2(new_n664), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n311), .B2(new_n351), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n311), .A2(new_n351), .A3(new_n1141), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n890), .B2(G330), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1072), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n880), .B1(new_n902), .B2(new_n903), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n1150), .C1(new_n1151), .C2(KEYINPUT40), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1139), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n890), .A2(G330), .A3(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1087), .A2(new_n904), .B1(new_n657), .B2(new_n664), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1088), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .A4(KEYINPUT120), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n727), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n731), .B1(G50), .B2(new_n807), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n756), .A2(new_n478), .B1(new_n766), .B2(new_n202), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G97), .B2(new_n757), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n459), .A2(new_n294), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G283), .B2(new_n979), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n779), .A2(G107), .B1(new_n809), .B2(new_n361), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n781), .A2(G68), .B1(new_n834), .B2(new_n784), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1166), .B(new_n246), .C1(G33), .C2(G41), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n757), .A2(G132), .B1(new_n809), .B2(G137), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT118), .Z(new_n1176));
  OAI22_X1  g0976(.A1(new_n770), .A2(new_n1120), .B1(new_n764), .B2(new_n1123), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT119), .Z(new_n1178));
  AOI22_X1  g0978(.A1(G150), .A2(new_n781), .B1(new_n755), .B2(G125), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n976), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n979), .C2(G124), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1174), .B1(new_n1171), .B2(new_n1170), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1163), .B1(new_n1186), .B2(new_n739), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1148), .B2(new_n736), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT121), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT121), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1162), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1160), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n920), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1094), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n693), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1094), .B1(new_n1092), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1194), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1193), .A2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1067), .A2(new_n735), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n731), .B1(G68), .B2(new_n807), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n756), .A2(new_n815), .B1(new_n764), .B2(new_n208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G77), .B2(new_n976), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n284), .B1(new_n979), .B2(G303), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n779), .A2(G283), .B1(new_n809), .B2(G107), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n361), .A2(new_n781), .B1(new_n757), .B2(G116), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT123), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n756), .A2(new_n826), .B1(new_n246), .B2(new_n761), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G159), .B2(new_n784), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n769), .A2(new_n254), .B1(new_n751), .B2(new_n1120), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n459), .B(new_n1219), .C1(G137), .C2(new_n779), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n757), .A2(new_n1124), .B1(new_n976), .B2(G58), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1216), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1208), .B1(new_n1224), .B2(new_n739), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT124), .Z(new_n1226));
  AOI22_X1  g1026(.A1(new_n1201), .A2(new_n727), .B1(new_n1207), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1097), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1228), .B(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1100), .A2(new_n955), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(G381));
  OR3_X1    g1032(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT125), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1110), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1107), .A2(KEYINPUT113), .A3(new_n1108), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1136), .B1(new_n1238), .B2(new_n1101), .ZN(new_n1239));
  INV_X1    g1039(.A(G375), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1235), .A2(new_n1239), .A3(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n665), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1239), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1193), .A2(new_n1205), .A3(G378), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1202), .A2(new_n1203), .A3(new_n955), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1188), .B1(new_n1249), .B2(new_n726), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1239), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1243), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(KEYINPUT126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT126), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1228), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n693), .B1(new_n1257), .B2(KEYINPUT60), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n1230), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1254), .B(new_n1256), .C1(new_n1260), .C2(new_n1227), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1253), .A4(new_n1227), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G2897), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1261), .A2(new_n1263), .B1(new_n1264), .B2(new_n1242), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1254), .B1(new_n1260), .B2(new_n1227), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1255), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(G2897), .A3(new_n1243), .A4(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1246), .B1(new_n1252), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1242), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1262), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1272), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G390), .B1(new_n971), .B2(new_n997), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n971), .A2(new_n997), .A3(G390), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(G396), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1278), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1279), .A2(new_n1283), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1271), .A2(new_n1277), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1252), .A2(new_n1290), .A3(new_n1275), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1252), .B2(new_n1275), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1291), .A2(new_n1270), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1293), .B2(new_n1287), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1239), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1247), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1285), .A2(new_n1275), .A3(new_n1286), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1275), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1287), .A2(new_n1276), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1296), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1285), .A2(new_n1275), .A3(new_n1286), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(G402));
endmodule


