

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764;

  NOR2_X1 U376 ( .A1(n635), .A2(n634), .ZN(n638) );
  XNOR2_X1 U377 ( .A(n379), .B(n477), .ZN(n597) );
  XNOR2_X1 U378 ( .A(n476), .B(n475), .ZN(n636) );
  NOR2_X1 U379 ( .A1(n531), .A2(n669), .ZN(n449) );
  XNOR2_X2 U380 ( .A(n503), .B(KEYINPUT4), .ZN(n511) );
  XNOR2_X1 U381 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n434) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n483) );
  XOR2_X1 U383 ( .A(KEYINPUT8), .B(n438), .Z(n500) );
  INV_X2 U384 ( .A(G953), .ZN(n755) );
  XOR2_X1 U385 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n354) );
  XOR2_X1 U386 ( .A(G116), .B(G101), .Z(n355) );
  XNOR2_X2 U387 ( .A(n582), .B(n581), .ZN(n645) );
  OR2_X2 U388 ( .A1(n608), .A2(n607), .ZN(n610) );
  NOR2_X1 U389 ( .A1(n599), .A2(n595), .ZN(n596) );
  NAND2_X1 U390 ( .A1(n656), .A2(n660), .ZN(n686) );
  OR2_X1 U391 ( .A1(n763), .A2(n600), .ZN(n601) );
  XNOR2_X1 U392 ( .A(n596), .B(KEYINPUT32), .ZN(n763) );
  OR2_X1 U393 ( .A1(n649), .A2(KEYINPUT44), .ZN(n600) );
  XNOR2_X1 U394 ( .A(n552), .B(n551), .ZN(n573) );
  XNOR2_X1 U395 ( .A(n524), .B(n523), .ZN(n656) );
  XNOR2_X1 U396 ( .A(n448), .B(n447), .ZN(n531) );
  AND2_X1 U397 ( .A1(n395), .A2(n358), .ZN(n396) );
  XNOR2_X1 U398 ( .A(n394), .B(n393), .ZN(n513) );
  XNOR2_X1 U399 ( .A(n355), .B(n470), .ZN(n394) );
  XNOR2_X1 U400 ( .A(n357), .B(n510), .ZN(n420) );
  XNOR2_X1 U401 ( .A(n392), .B(G104), .ZN(n514) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(G113), .ZN(n470) );
  BUF_X1 U403 ( .A(n525), .Z(n356) );
  XNOR2_X1 U404 ( .A(n521), .B(KEYINPUT39), .ZN(n525) );
  NAND2_X1 U405 ( .A1(n525), .A2(n654), .ZN(n527) );
  XNOR2_X1 U406 ( .A(n511), .B(n458), .ZN(n476) );
  INV_X1 U407 ( .A(G134), .ZN(n457) );
  XNOR2_X1 U408 ( .A(n513), .B(n389), .ZN(n738) );
  XNOR2_X1 U409 ( .A(n514), .B(n390), .ZN(n389) );
  XNOR2_X1 U410 ( .A(n391), .B(KEYINPUT16), .ZN(n390) );
  XNOR2_X1 U411 ( .A(KEYINPUT70), .B(G122), .ZN(n391) );
  XNOR2_X1 U412 ( .A(n563), .B(KEYINPUT38), .ZN(n680) );
  NAND2_X1 U413 ( .A1(n418), .A2(n417), .ZN(n552) );
  INV_X1 U414 ( .A(n563), .ZN(n418) );
  NAND2_X1 U415 ( .A1(n376), .A2(n373), .ZN(n528) );
  OR2_X1 U416 ( .A1(n725), .A2(n374), .ZN(n373) );
  AND2_X1 U417 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U418 ( .A1(n494), .A2(n375), .ZN(n374) );
  NAND2_X1 U419 ( .A1(G472), .A2(n375), .ZN(n398) );
  XNOR2_X1 U420 ( .A(n421), .B(n420), .ZN(n512) );
  XNOR2_X1 U421 ( .A(n509), .B(n354), .ZN(n421) );
  NOR2_X1 U422 ( .A1(n412), .A2(n611), .ZN(n411) );
  NOR2_X1 U423 ( .A1(n558), .A2(n381), .ZN(n380) );
  NAND2_X1 U424 ( .A1(n662), .A2(n557), .ZN(n381) );
  NAND2_X1 U425 ( .A1(n725), .A2(n424), .ZN(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT101), .B(KEYINPUT98), .Z(n489) );
  XNOR2_X1 U427 ( .A(G131), .B(G140), .ZN(n488) );
  XNOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n366) );
  XOR2_X1 U429 ( .A(G122), .B(G104), .Z(n487) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n516) );
  XNOR2_X1 U431 ( .A(n574), .B(KEYINPUT0), .ZN(n589) );
  NOR2_X1 U432 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U433 ( .A1(n444), .A2(n375), .ZN(n448) );
  XNOR2_X1 U434 ( .A(G137), .B(G146), .ZN(n472) );
  XNOR2_X1 U435 ( .A(n440), .B(n409), .ZN(n408) );
  INV_X1 U436 ( .A(KEYINPUT93), .ZN(n409) );
  XNOR2_X1 U437 ( .A(G119), .B(G110), .ZN(n442) );
  XNOR2_X1 U438 ( .A(n429), .B(G902), .ZN(n633) );
  INV_X1 U439 ( .A(KEYINPUT15), .ZN(n429) );
  INV_X1 U440 ( .A(KEYINPUT72), .ZN(n568) );
  XNOR2_X1 U441 ( .A(G110), .B(G107), .ZN(n392) );
  XNOR2_X1 U442 ( .A(n476), .B(n459), .ZN(n752) );
  XNOR2_X1 U443 ( .A(n388), .B(n530), .ZN(n699) );
  INV_X1 U444 ( .A(KEYINPUT41), .ZN(n530) );
  NAND2_X1 U445 ( .A1(n680), .A2(n387), .ZN(n388) );
  AND2_X1 U446 ( .A1(n481), .A2(n680), .ZN(n427) );
  INV_X1 U447 ( .A(n666), .ZN(n425) );
  NAND2_X1 U448 ( .A1(n552), .A2(KEYINPUT36), .ZN(n370) );
  NOR2_X1 U449 ( .A1(n560), .A2(n372), .ZN(n371) );
  OR2_X1 U450 ( .A1(n552), .A2(KEYINPUT36), .ZN(n372) );
  XOR2_X1 U451 ( .A(n628), .B(n627), .Z(n629) );
  XNOR2_X1 U452 ( .A(n539), .B(KEYINPUT64), .ZN(n540) );
  XNOR2_X1 U453 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n365) );
  NAND2_X1 U454 ( .A1(n424), .A2(G902), .ZN(n377) );
  XNOR2_X1 U455 ( .A(n469), .B(KEYINPUT87), .ZN(n393) );
  XNOR2_X1 U456 ( .A(KEYINPUT69), .B(G119), .ZN(n469) );
  XNOR2_X1 U457 ( .A(G128), .B(KEYINPUT23), .ZN(n435) );
  AND2_X1 U458 ( .A1(n680), .A2(n417), .ZN(n687) );
  NAND2_X1 U459 ( .A1(G234), .A2(G237), .ZN(n450) );
  OR2_X1 U460 ( .A1(n602), .A2(n665), .ZN(n603) );
  INV_X1 U461 ( .A(n362), .ZN(n576) );
  XNOR2_X1 U462 ( .A(G107), .B(KEYINPUT9), .ZN(n496) );
  XOR2_X1 U463 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n497) );
  XNOR2_X1 U464 ( .A(G116), .B(G134), .ZN(n495) );
  XNOR2_X1 U465 ( .A(n493), .B(n492), .ZN(n725) );
  BUF_X1 U466 ( .A(n589), .Z(n605) );
  XNOR2_X1 U467 ( .A(n517), .B(KEYINPUT75), .ZN(n518) );
  XNOR2_X1 U468 ( .A(n528), .B(n423), .ZN(n522) );
  INV_X1 U469 ( .A(KEYINPUT102), .ZN(n423) );
  XNOR2_X1 U470 ( .A(n419), .B(n359), .ZN(n593) );
  AND2_X1 U471 ( .A1(n684), .A2(n587), .ZN(n588) );
  BUF_X1 U472 ( .A(n531), .Z(n668) );
  XNOR2_X1 U473 ( .A(n433), .B(n439), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n408), .B(n443), .ZN(n407) );
  XNOR2_X1 U475 ( .A(KEYINPUT91), .B(G101), .ZN(n461) );
  XNOR2_X1 U476 ( .A(n538), .B(n384), .ZN(n764) );
  NOR2_X1 U477 ( .A1(n699), .A2(n553), .ZN(n538) );
  NAND2_X1 U478 ( .A1(n368), .A2(n367), .ZN(n662) );
  NOR2_X1 U479 ( .A1(n371), .A2(n369), .ZN(n368) );
  NAND2_X1 U480 ( .A1(n425), .A2(n370), .ZN(n369) );
  INV_X1 U481 ( .A(KEYINPUT60), .ZN(n399) );
  NAND2_X1 U482 ( .A1(n401), .A2(n404), .ZN(n400) );
  XNOR2_X1 U483 ( .A(n402), .B(n728), .ZN(n401) );
  NAND2_X1 U484 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U485 ( .A(n406), .B(n629), .ZN(n405) );
  XNOR2_X1 U486 ( .A(n478), .B(KEYINPUT89), .ZN(n682) );
  INV_X1 U487 ( .A(n682), .ZN(n417) );
  INV_X1 U488 ( .A(n494), .ZN(n424) );
  INV_X1 U489 ( .A(G902), .ZN(n375) );
  XOR2_X1 U490 ( .A(KEYINPUT88), .B(KEYINPUT74), .Z(n357) );
  NAND2_X1 U491 ( .A1(n634), .A2(G902), .ZN(n358) );
  XOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n359) );
  XOR2_X1 U493 ( .A(n479), .B(KEYINPUT109), .Z(n360) );
  INV_X1 U494 ( .A(n444), .ZN(n734) );
  XNOR2_X1 U495 ( .A(n407), .B(n410), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n361) );
  AND2_X1 U497 ( .A1(n630), .A2(G953), .ZN(n737) );
  INV_X1 U498 ( .A(n737), .ZN(n404) );
  XNOR2_X1 U499 ( .A(n363), .B(n466), .ZN(n362) );
  NOR2_X1 U500 ( .A1(n717), .A2(G902), .ZN(n363) );
  XNOR2_X1 U501 ( .A(n513), .B(n474), .ZN(n475) );
  XNOR2_X1 U502 ( .A(n515), .B(n738), .ZN(n628) );
  NOR2_X1 U503 ( .A1(n628), .A2(n633), .ZN(n519) );
  NAND2_X1 U504 ( .A1(n396), .A2(n397), .ZN(n364) );
  NAND2_X1 U505 ( .A1(n396), .A2(n397), .ZN(n379) );
  OR2_X1 U506 ( .A1(n636), .A2(n398), .ZN(n397) );
  XNOR2_X1 U507 ( .A(n366), .B(n365), .ZN(n386) );
  NAND2_X1 U508 ( .A1(n560), .A2(KEYINPUT36), .ZN(n367) );
  INV_X1 U509 ( .A(n364), .ZN(n579) );
  XNOR2_X1 U510 ( .A(n364), .B(KEYINPUT6), .ZN(n594) );
  OR2_X1 U511 ( .A1(n665), .A2(n364), .ZN(n583) );
  NAND2_X1 U512 ( .A1(n671), .A2(n364), .ZN(n672) );
  NAND2_X1 U513 ( .A1(n382), .A2(n380), .ZN(n385) );
  XNOR2_X1 U514 ( .A(n383), .B(n540), .ZN(n382) );
  NAND2_X1 U515 ( .A1(n632), .A2(n764), .ZN(n383) );
  INV_X1 U516 ( .A(KEYINPUT42), .ZN(n384) );
  XNOR2_X2 U517 ( .A(n527), .B(n526), .ZN(n632) );
  XNOR2_X1 U518 ( .A(n752), .B(n464), .ZN(n717) );
  INV_X1 U519 ( .A(G140), .ZN(n441) );
  XNOR2_X1 U520 ( .A(n386), .B(n422), .ZN(n485) );
  XNOR2_X1 U521 ( .A(n385), .B(n559), .ZN(n565) );
  XNOR2_X1 U522 ( .A(n480), .B(n360), .ZN(n481) );
  NOR2_X1 U523 ( .A1(n656), .A2(n602), .ZN(n547) );
  NAND2_X2 U524 ( .A1(n625), .A2(n707), .ZN(n724) );
  NAND2_X1 U525 ( .A1(n697), .A2(n605), .ZN(n606) );
  XNOR2_X2 U526 ( .A(n604), .B(KEYINPUT33), .ZN(n697) );
  XNOR2_X2 U527 ( .A(n576), .B(KEYINPUT1), .ZN(n666) );
  AND2_X1 U528 ( .A1(n684), .A2(n417), .ZN(n387) );
  NAND2_X1 U529 ( .A1(n636), .A2(n634), .ZN(n395) );
  XNOR2_X1 U530 ( .A(n400), .B(n399), .ZN(G60) );
  NAND2_X1 U531 ( .A1(n724), .A2(n723), .ZN(n402) );
  XNOR2_X1 U532 ( .A(n403), .B(n361), .ZN(G51) );
  NAND2_X1 U533 ( .A1(n729), .A2(G210), .ZN(n406) );
  NAND2_X1 U534 ( .A1(n414), .A2(n411), .ZN(n618) );
  AND2_X1 U535 ( .A1(n413), .A2(n631), .ZN(n412) );
  XNOR2_X2 U536 ( .A(n610), .B(n609), .ZN(n631) );
  NAND2_X1 U537 ( .A1(n601), .A2(KEYINPUT84), .ZN(n413) );
  NAND2_X1 U538 ( .A1(n415), .A2(n616), .ZN(n414) );
  NAND2_X1 U539 ( .A1(n416), .A2(n614), .ZN(n415) );
  NAND2_X1 U540 ( .A1(n612), .A2(KEYINPUT84), .ZN(n416) );
  XNOR2_X2 U541 ( .A(n519), .B(n518), .ZN(n563) );
  NAND2_X1 U542 ( .A1(n593), .A2(n668), .ZN(n599) );
  NAND2_X1 U543 ( .A1(n589), .A2(n588), .ZN(n419) );
  NAND2_X1 U544 ( .A1(n483), .A2(G214), .ZN(n422) );
  XNOR2_X2 U545 ( .A(n426), .B(n456), .ZN(n503) );
  XNOR2_X2 U546 ( .A(G143), .B(KEYINPUT65), .ZN(n426) );
  NAND2_X1 U547 ( .A1(n427), .A2(n482), .ZN(n521) );
  AND2_X1 U548 ( .A1(n481), .A2(n482), .ZN(n428) );
  NAND2_X1 U549 ( .A1(n428), .A2(n520), .ZN(n541) );
  BUF_X1 U550 ( .A(n706), .Z(n754) );
  INV_X1 U551 ( .A(n680), .ZN(n681) );
  INV_X1 U552 ( .A(n437), .ZN(n440) );
  XNOR2_X1 U553 ( .A(n485), .B(n750), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n432) );
  INV_X1 U555 ( .A(n633), .ZN(n722) );
  NAND2_X1 U556 ( .A1(G234), .A2(n722), .ZN(n430) );
  XNOR2_X1 U557 ( .A(KEYINPUT20), .B(n430), .ZN(n445) );
  NAND2_X1 U558 ( .A1(n445), .A2(G221), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n432), .B(n431), .ZN(n669) );
  XNOR2_X2 U560 ( .A(G146), .B(G125), .ZN(n508) );
  XNOR2_X1 U561 ( .A(n508), .B(KEYINPUT10), .ZN(n484) );
  XNOR2_X1 U562 ( .A(n484), .B(KEYINPUT24), .ZN(n433) );
  INV_X1 U563 ( .A(n434), .ZN(n436) );
  XNOR2_X1 U564 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U565 ( .A1(G234), .A2(n755), .ZN(n438) );
  NAND2_X1 U566 ( .A1(G221), .A2(n500), .ZN(n439) );
  XNOR2_X1 U567 ( .A(n441), .B(G137), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n442), .B(n459), .ZN(n443) );
  NAND2_X1 U569 ( .A1(n445), .A2(G217), .ZN(n446) );
  XNOR2_X1 U570 ( .A(n446), .B(KEYINPUT25), .ZN(n447) );
  XNOR2_X1 U571 ( .A(n449), .B(KEYINPUT67), .ZN(n575) );
  XNOR2_X1 U572 ( .A(n450), .B(KEYINPUT90), .ZN(n451) );
  XNOR2_X1 U573 ( .A(KEYINPUT14), .B(n451), .ZN(n454) );
  AND2_X1 U574 ( .A1(n454), .A2(G953), .ZN(n452) );
  NAND2_X1 U575 ( .A1(G902), .A2(n452), .ZN(n569) );
  XOR2_X1 U576 ( .A(n569), .B(KEYINPUT107), .Z(n453) );
  NOR2_X1 U577 ( .A1(n453), .A2(G900), .ZN(n455) );
  NAND2_X1 U578 ( .A1(G952), .A2(n454), .ZN(n696) );
  NOR2_X1 U579 ( .A1(n696), .A2(G953), .ZN(n570) );
  NOR2_X1 U580 ( .A1(n455), .A2(n570), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n575), .A2(n532), .ZN(n467) );
  INV_X1 U582 ( .A(G128), .ZN(n456) );
  XNOR2_X1 U583 ( .A(n457), .B(G131), .ZN(n458) );
  NAND2_X1 U584 ( .A1(n755), .A2(G227), .ZN(n460) );
  XNOR2_X1 U585 ( .A(n460), .B(G146), .ZN(n462) );
  XNOR2_X1 U586 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U587 ( .A(n514), .B(n463), .ZN(n464) );
  INV_X1 U588 ( .A(KEYINPUT68), .ZN(n465) );
  XNOR2_X1 U589 ( .A(n465), .B(G469), .ZN(n466) );
  NAND2_X1 U590 ( .A1(n467), .A2(n362), .ZN(n468) );
  XNOR2_X1 U591 ( .A(n468), .B(KEYINPUT73), .ZN(n482) );
  NAND2_X1 U592 ( .A1(n483), .A2(G210), .ZN(n471) );
  XNOR2_X1 U593 ( .A(n471), .B(KEYINPUT5), .ZN(n473) );
  XNOR2_X1 U594 ( .A(n473), .B(n472), .ZN(n474) );
  INV_X1 U595 ( .A(G472), .ZN(n634) );
  INV_X1 U596 ( .A(KEYINPUT105), .ZN(n477) );
  NAND2_X1 U597 ( .A1(G214), .A2(n516), .ZN(n478) );
  NOR2_X1 U598 ( .A1(n597), .A2(n682), .ZN(n480) );
  XNOR2_X1 U599 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n479) );
  BUF_X1 U600 ( .A(n484), .Z(n750) );
  XNOR2_X1 U601 ( .A(G113), .B(G143), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n487), .B(n486), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U604 ( .A(n491), .B(n490), .Z(n492) );
  XNOR2_X1 U605 ( .A(KEYINPUT13), .B(G475), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n495), .B(G122), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U608 ( .A(n499), .B(n498), .Z(n502) );
  NAND2_X1 U609 ( .A1(G217), .A2(n500), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n502), .B(n501), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n503), .B(n504), .ZN(n731) );
  NAND2_X1 U612 ( .A1(n731), .A2(n375), .ZN(n505) );
  XNOR2_X1 U613 ( .A(n505), .B(G478), .ZN(n529) );
  AND2_X1 U614 ( .A1(n528), .A2(n529), .ZN(n507) );
  INV_X1 U615 ( .A(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U616 ( .A(n507), .B(n506), .ZN(n607) );
  INV_X1 U617 ( .A(n508), .ZN(n509) );
  NAND2_X1 U618 ( .A1(G224), .A2(n755), .ZN(n510) );
  XNOR2_X1 U619 ( .A(n511), .B(n512), .ZN(n515) );
  NAND2_X1 U620 ( .A1(G210), .A2(n516), .ZN(n517) );
  NOR2_X1 U621 ( .A1(n607), .A2(n563), .ZN(n520) );
  XNOR2_X1 U622 ( .A(n541), .B(G143), .ZN(G45) );
  NAND2_X1 U623 ( .A1(n522), .A2(n529), .ZN(n660) );
  INV_X1 U624 ( .A(n660), .ZN(n650) );
  NAND2_X1 U625 ( .A1(n356), .A2(n650), .ZN(n620) );
  XNOR2_X1 U626 ( .A(n620), .B(G134), .ZN(G36) );
  NOR2_X1 U627 ( .A1(n522), .A2(n529), .ZN(n524) );
  INV_X1 U628 ( .A(KEYINPUT104), .ZN(n523) );
  INV_X1 U629 ( .A(n656), .ZN(n654) );
  XOR2_X1 U630 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n526) );
  NOR2_X1 U631 ( .A1(n529), .A2(n528), .ZN(n684) );
  NOR2_X1 U632 ( .A1(n532), .A2(n669), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n668), .A2(n533), .ZN(n545) );
  NOR2_X1 U634 ( .A1(n597), .A2(n545), .ZN(n535) );
  XNOR2_X1 U635 ( .A(KEYINPUT112), .B(KEYINPUT28), .ZN(n534) );
  XNOR2_X1 U636 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n576), .B(KEYINPUT111), .ZN(n536) );
  NAND2_X1 U638 ( .A1(n537), .A2(n536), .ZN(n553) );
  XNOR2_X1 U639 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n541), .B(KEYINPUT78), .ZN(n543) );
  INV_X1 U641 ( .A(n686), .ZN(n549) );
  NAND2_X1 U642 ( .A1(n549), .A2(KEYINPUT47), .ZN(n542) );
  NAND2_X1 U643 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U644 ( .A(KEYINPUT76), .B(n544), .ZN(n558) );
  INV_X1 U645 ( .A(n594), .ZN(n602) );
  INV_X1 U646 ( .A(n545), .ZN(n546) );
  NAND2_X1 U647 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U648 ( .A(n548), .B(KEYINPUT108), .ZN(n560) );
  NOR2_X1 U649 ( .A1(KEYINPUT47), .A2(n549), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT71), .ZN(n554) );
  INV_X1 U651 ( .A(KEYINPUT19), .ZN(n551) );
  NOR2_X1 U652 ( .A1(n553), .A2(n573), .ZN(n653) );
  NAND2_X1 U653 ( .A1(n554), .A2(n653), .ZN(n556) );
  OR2_X1 U654 ( .A1(KEYINPUT47), .A2(n653), .ZN(n555) );
  NAND2_X1 U655 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U656 ( .A(KEYINPUT48), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n560), .A2(n682), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n561), .A2(n666), .ZN(n562) );
  XNOR2_X1 U659 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  NAND2_X1 U660 ( .A1(n564), .A2(n563), .ZN(n664) );
  NAND2_X1 U661 ( .A1(n565), .A2(n664), .ZN(n566) );
  XNOR2_X1 U662 ( .A(n566), .B(KEYINPUT81), .ZN(n621) );
  NAND2_X1 U663 ( .A1(n621), .A2(n620), .ZN(n567) );
  XNOR2_X2 U664 ( .A(n567), .B(KEYINPUT80), .ZN(n706) );
  XNOR2_X1 U665 ( .A(n706), .B(n568), .ZN(n619) );
  NOR2_X1 U666 ( .A1(G898), .A2(n569), .ZN(n571) );
  NOR2_X1 U667 ( .A1(n571), .A2(n570), .ZN(n572) );
  BUF_X1 U668 ( .A(n575), .Z(n665) );
  NOR2_X1 U669 ( .A1(n576), .A2(n665), .ZN(n577) );
  NAND2_X1 U670 ( .A1(n605), .A2(n577), .ZN(n578) );
  XNOR2_X1 U671 ( .A(n578), .B(KEYINPUT96), .ZN(n580) );
  OR2_X1 U672 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U673 ( .A(KEYINPUT97), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n666), .A2(n583), .ZN(n675) );
  NAND2_X1 U675 ( .A1(n605), .A2(n675), .ZN(n585) );
  INV_X1 U676 ( .A(KEYINPUT31), .ZN(n584) );
  XNOR2_X1 U677 ( .A(n585), .B(n584), .ZN(n659) );
  NAND2_X1 U678 ( .A1(n645), .A2(n659), .ZN(n586) );
  NAND2_X1 U679 ( .A1(n586), .A2(n686), .ZN(n592) );
  INV_X1 U680 ( .A(n669), .ZN(n587) );
  NOR2_X1 U681 ( .A1(n594), .A2(n668), .ZN(n590) );
  AND2_X1 U682 ( .A1(n666), .A2(n590), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n593), .A2(n591), .ZN(n642) );
  NAND2_X1 U684 ( .A1(n592), .A2(n642), .ZN(n611) );
  OR2_X1 U685 ( .A1(n666), .A2(n594), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n666), .A2(n597), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n649) );
  OR2_X1 U688 ( .A1(n666), .A2(n603), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n606), .B(KEYINPUT34), .ZN(n608) );
  INV_X1 U690 ( .A(KEYINPUT35), .ZN(n609) );
  INV_X1 U691 ( .A(n631), .ZN(n612) );
  INV_X1 U692 ( .A(KEYINPUT44), .ZN(n615) );
  OR2_X1 U693 ( .A1(n649), .A2(n615), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n763), .A2(n613), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(KEYINPUT84), .ZN(n616) );
  INV_X1 U696 ( .A(KEYINPUT45), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n618), .B(n617), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n622), .A2(KEYINPUT2), .ZN(n704) );
  NAND2_X1 U699 ( .A1(n619), .A2(n704), .ZN(n625) );
  AND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n623) );
  INV_X1 U701 ( .A(n622), .ZN(n741) );
  NAND2_X1 U702 ( .A1(n623), .A2(n741), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n624), .A2(KEYINPUT2), .ZN(n707) );
  AND2_X2 U704 ( .A1(n724), .A2(n633), .ZN(n729) );
  XNOR2_X1 U705 ( .A(KEYINPUT77), .B(KEYINPUT54), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT55), .ZN(n627) );
  INV_X1 U707 ( .A(G952), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n631), .B(G122), .ZN(G24) );
  XNOR2_X1 U709 ( .A(n632), .B(G131), .ZN(G33) );
  NAND2_X1 U710 ( .A1(n724), .A2(n633), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT62), .B(n636), .Z(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n639), .A2(n737), .ZN(n641) );
  XNOR2_X1 U714 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(G57) );
  XNOR2_X1 U716 ( .A(G101), .B(KEYINPUT114), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(G3) );
  NOR2_X1 U718 ( .A1(n656), .A2(n645), .ZN(n644) );
  XOR2_X1 U719 ( .A(G104), .B(n644), .Z(G6) );
  NOR2_X1 U720 ( .A1(n660), .A2(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U723 ( .A(G107), .B(n648), .ZN(G9) );
  XOR2_X1 U724 ( .A(G110), .B(n649), .Z(G12) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .Z(n652) );
  NAND2_X1 U726 ( .A1(n653), .A2(n650), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(G30) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(G146), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n656), .A2(n659), .ZN(n658) );
  XNOR2_X1 U731 ( .A(G113), .B(KEYINPUT115), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(G15) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U734 ( .A(G116), .B(n661), .Z(G18) );
  XOR2_X1 U735 ( .A(n662), .B(G125), .Z(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U737 ( .A(G140), .B(n664), .ZN(G42) );
  XOR2_X1 U738 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n694) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT50), .B(n667), .Z(n673) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT49), .B(n670), .Z(n671) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT116), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n677), .Z(n678) );
  NOR2_X1 U747 ( .A1(n699), .A2(n678), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(KEYINPUT117), .ZN(n692) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT118), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n690), .A2(n697), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U756 ( .A(n694), .B(n693), .Z(n695) );
  NOR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U758 ( .A(n697), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U761 ( .A(n702), .B(KEYINPUT120), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n703), .A2(n755), .ZN(n713) );
  NOR2_X1 U763 ( .A1(n704), .A2(KEYINPUT2), .ZN(n705) );
  XOR2_X1 U764 ( .A(KEYINPUT79), .B(n705), .Z(n711) );
  NOR2_X1 U765 ( .A1(n754), .A2(KEYINPUT2), .ZN(n709) );
  INV_X1 U766 ( .A(n707), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U770 ( .A(KEYINPUT53), .B(n714), .ZN(G75) );
  BUF_X1 U771 ( .A(n729), .Z(n733) );
  NAND2_X1 U772 ( .A1(n733), .A2(G469), .ZN(n719) );
  XOR2_X1 U773 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XOR2_X1 U774 ( .A(n715), .B(KEYINPUT121), .Z(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U776 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n737), .A2(n720), .ZN(G54) );
  INV_X1 U778 ( .A(G475), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U780 ( .A(KEYINPUT59), .B(KEYINPUT86), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT122), .ZN(n726) );
  XNOR2_X1 U782 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U783 ( .A1(n729), .A2(G478), .ZN(n730) );
  XOR2_X1 U784 ( .A(n731), .B(n730), .Z(n732) );
  NOR2_X1 U785 ( .A1(n737), .A2(n732), .ZN(G63) );
  NAND2_X1 U786 ( .A1(n733), .A2(G217), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U788 ( .A1(n737), .A2(n736), .ZN(G66) );
  NOR2_X1 U789 ( .A1(G898), .A2(n755), .ZN(n740) );
  XOR2_X1 U790 ( .A(n738), .B(KEYINPUT124), .Z(n739) );
  NOR2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n749) );
  BUF_X1 U792 ( .A(n741), .Z(n742) );
  NAND2_X1 U793 ( .A1(n742), .A2(n755), .ZN(n747) );
  XOR2_X1 U794 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n744) );
  NAND2_X1 U795 ( .A1(G224), .A2(G953), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U798 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U799 ( .A(n749), .B(n748), .ZN(G69) );
  XNOR2_X1 U800 ( .A(n750), .B(KEYINPUT125), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n757) );
  XNOR2_X1 U802 ( .A(n757), .B(KEYINPUT126), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n761) );
  XNOR2_X1 U805 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U809 ( .A(KEYINPUT127), .B(n762), .Z(G72) );
  XOR2_X1 U810 ( .A(n763), .B(G119), .Z(G21) );
  XNOR2_X1 U811 ( .A(G137), .B(n764), .ZN(G39) );
endmodule

