

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739;

  NAND2_X1 U361 ( .A1(n433), .A2(n436), .ZN(n662) );
  XNOR2_X1 U362 ( .A(n348), .B(G128), .ZN(n503) );
  XNOR2_X2 U363 ( .A(n468), .B(n467), .ZN(n543) );
  XNOR2_X2 U364 ( .A(n555), .B(KEYINPUT33), .ZN(n686) );
  AND2_X2 U365 ( .A1(n362), .A2(n654), .ZN(n555) );
  XNOR2_X2 U366 ( .A(G110), .B(G104), .ZN(n482) );
  XNOR2_X2 U367 ( .A(n592), .B(KEYINPUT1), .ZN(n654) );
  XNOR2_X2 U368 ( .A(n391), .B(n509), .ZN(n593) );
  XNOR2_X1 U369 ( .A(n376), .B(n402), .ZN(n375) );
  NOR2_X1 U370 ( .A1(n624), .A2(n709), .ZN(n625) );
  NOR2_X1 U371 ( .A1(n703), .A2(n709), .ZN(n407) );
  NOR2_X1 U372 ( .A1(n696), .A2(n709), .ZN(n698) );
  NAND2_X1 U373 ( .A1(n418), .A2(n622), .ZN(n417) );
  NAND2_X1 U374 ( .A1(n728), .A2(n449), .ZN(n418) );
  NAND2_X1 U375 ( .A1(n375), .A2(n409), .ZN(n728) );
  NOR2_X1 U376 ( .A1(n601), .A2(n398), .ZN(n602) );
  INV_X1 U377 ( .A(n651), .ZN(n410) );
  INV_X1 U378 ( .A(G902), .ZN(n343) );
  INV_X1 U379 ( .A(G143), .ZN(n348) );
  NOR2_X1 U380 ( .A1(n410), .A2(n738), .ZN(n409) );
  AND2_X1 U381 ( .A1(n372), .A2(n565), .ZN(n566) );
  XNOR2_X1 U382 ( .A(n419), .B(n358), .ZN(n608) );
  XNOR2_X1 U383 ( .A(n544), .B(KEYINPUT68), .ZN(n655) );
  NAND2_X1 U384 ( .A1(n585), .A2(n671), .ZN(n445) );
  NAND2_X2 U385 ( .A1(n344), .A2(n341), .ZN(n592) );
  AND2_X1 U386 ( .A1(n346), .A2(n345), .ZN(n344) );
  XNOR2_X1 U387 ( .A(n504), .B(n393), .ZN(n447) );
  XNOR2_X1 U388 ( .A(n500), .B(n394), .ZN(n393) );
  NAND2_X1 U389 ( .A1(n489), .A2(n343), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n503), .B(G134), .ZN(n373) );
  NAND2_X1 U391 ( .A1(n347), .A2(G902), .ZN(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT69), .B(G131), .Z(n486) );
  XNOR2_X2 U393 ( .A(n340), .B(n516), .ZN(n556) );
  NOR2_X2 U394 ( .A1(n593), .A2(n515), .ZN(n340) );
  XNOR2_X2 U395 ( .A(n445), .B(KEYINPUT86), .ZN(n391) );
  NOR2_X2 U396 ( .A1(n365), .A2(n636), .ZN(n567) );
  XNOR2_X2 U397 ( .A(n367), .B(n385), .ZN(n365) );
  OR2_X1 U398 ( .A1(n700), .A2(n342), .ZN(n341) );
  NAND2_X1 U399 ( .A1(n700), .A2(n347), .ZN(n346) );
  INV_X1 U400 ( .A(n489), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n403), .B(n488), .ZN(n700) );
  NOR2_X1 U402 ( .A1(n443), .A2(n417), .ZN(n349) );
  BUF_X1 U403 ( .A(n693), .Z(n350) );
  NOR2_X1 U404 ( .A1(n443), .A2(n417), .ZN(n416) );
  XNOR2_X1 U405 ( .A(n447), .B(n446), .ZN(n693) );
  AND2_X1 U406 ( .A1(n416), .A2(n441), .ZN(n363) );
  XNOR2_X1 U407 ( .A(n395), .B(G125), .ZN(n497) );
  INV_X1 U408 ( .A(G146), .ZN(n395) );
  AND2_X1 U409 ( .A1(n374), .A2(n437), .ZN(n436) );
  NAND2_X1 U410 ( .A1(G472), .A2(G902), .ZN(n437) );
  NAND2_X1 U411 ( .A1(n444), .A2(n435), .ZN(n434) );
  INV_X1 U412 ( .A(G902), .ZN(n435) );
  INV_X1 U413 ( .A(n486), .ZN(n390) );
  XNOR2_X1 U414 ( .A(n727), .B(G101), .ZN(n491) );
  NOR2_X1 U415 ( .A1(n590), .A2(n589), .ZN(n613) );
  NOR2_X1 U416 ( .A1(n543), .A2(n590), .ZN(n544) );
  XNOR2_X1 U417 ( .A(G122), .B(KEYINPUT9), .ZN(n524) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n492) );
  XNOR2_X1 U419 ( .A(G113), .B(G122), .ZN(n474) );
  XOR2_X1 U420 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n475) );
  XNOR2_X1 U421 ( .A(KEYINPUT10), .B(G140), .ZN(n472) );
  XNOR2_X1 U422 ( .A(G137), .B(KEYINPUT70), .ZN(n532) );
  INV_X1 U423 ( .A(KEYINPUT73), .ZN(n568) );
  NAND2_X1 U424 ( .A1(n428), .A2(n425), .ZN(n581) );
  AND2_X1 U425 ( .A1(n431), .A2(n355), .ZN(n428) );
  OR2_X1 U426 ( .A1(n705), .A2(G902), .ZN(n467) );
  INV_X1 U427 ( .A(KEYINPUT96), .ZN(n469) );
  XNOR2_X1 U428 ( .A(KEYINPUT0), .B(KEYINPUT87), .ZN(n516) );
  XNOR2_X1 U429 ( .A(n424), .B(n422), .ZN(n494) );
  XNOR2_X1 U430 ( .A(n354), .B(n423), .ZN(n422) );
  XNOR2_X1 U431 ( .A(n502), .B(n491), .ZN(n424) );
  XNOR2_X1 U432 ( .A(n461), .B(n460), .ZN(n459) );
  XNOR2_X1 U433 ( .A(G128), .B(G119), .ZN(n460) );
  XNOR2_X1 U434 ( .A(n462), .B(G110), .ZN(n461) );
  INV_X1 U435 ( .A(KEYINPUT24), .ZN(n462) );
  XNOR2_X1 U436 ( .A(n458), .B(n457), .ZN(n456) );
  XNOR2_X1 U437 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U438 ( .A(KEYINPUT77), .B(KEYINPUT23), .ZN(n457) );
  XNOR2_X1 U439 ( .A(n528), .B(n413), .ZN(n704) );
  XNOR2_X1 U440 ( .A(G116), .B(G107), .ZN(n526) );
  XNOR2_X1 U441 ( .A(n725), .B(G146), .ZN(n495) );
  INV_X1 U442 ( .A(G140), .ZN(n487) );
  NAND2_X1 U443 ( .A1(n596), .A2(n672), .ZN(n419) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n387) );
  INV_X1 U445 ( .A(KEYINPUT106), .ZN(n388) );
  OR2_X1 U446 ( .A1(n616), .A2(n658), .ZN(n389) );
  NAND2_X1 U447 ( .A1(n654), .A2(n655), .ZN(n553) );
  INV_X1 U448 ( .A(KEYINPUT83), .ZN(n399) );
  NAND2_X1 U449 ( .A1(n671), .A2(n430), .ZN(n429) );
  XNOR2_X1 U450 ( .A(n519), .B(n518), .ZN(n538) );
  XOR2_X1 U451 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n519) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n517) );
  INV_X1 U453 ( .A(KEYINPUT15), .ZN(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT89), .B(G902), .ZN(n401) );
  INV_X1 U455 ( .A(KEYINPUT30), .ZN(n430) );
  AND2_X1 U456 ( .A1(n433), .A2(KEYINPUT30), .ZN(n432) );
  XNOR2_X1 U457 ( .A(n493), .B(G137), .ZN(n423) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n727) );
  XNOR2_X1 U459 ( .A(n353), .B(n490), .ZN(n502) );
  XNOR2_X1 U460 ( .A(G119), .B(KEYINPUT3), .ZN(n490) );
  XNOR2_X1 U461 ( .A(n525), .B(n411), .ZN(n527) );
  XNOR2_X1 U462 ( .A(n524), .B(n412), .ZN(n411) );
  INV_X1 U463 ( .A(KEYINPUT7), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n396), .B(n497), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n496), .B(KEYINPUT80), .ZN(n396) );
  NAND2_X1 U466 ( .A1(G224), .A2(n729), .ZN(n496) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n498) );
  XOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n499) );
  NAND2_X1 U469 ( .A1(n378), .A2(n377), .ZN(n376) );
  AND2_X1 U470 ( .A1(n421), .A2(n612), .ZN(n378) );
  XNOR2_X1 U471 ( .A(n609), .B(KEYINPUT46), .ZN(n610) );
  INV_X1 U472 ( .A(KEYINPUT48), .ZN(n402) );
  NOR2_X1 U473 ( .A1(G902), .A2(G237), .ZN(n505) );
  XNOR2_X1 U474 ( .A(n502), .B(n501), .ZN(n716) );
  XNOR2_X1 U475 ( .A(KEYINPUT16), .B(G122), .ZN(n501) );
  NAND2_X1 U476 ( .A1(n448), .A2(n442), .ZN(n441) );
  NOR2_X1 U477 ( .A1(n728), .A2(n449), .ZN(n448) );
  XNOR2_X1 U478 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U479 ( .A(n476), .B(n470), .ZN(n477) );
  NAND2_X1 U480 ( .A1(G214), .A2(n508), .ZN(n671) );
  XNOR2_X1 U481 ( .A(n646), .B(n408), .ZN(n586) );
  INV_X1 U482 ( .A(KEYINPUT103), .ZN(n408) );
  XNOR2_X1 U483 ( .A(n654), .B(n454), .ZN(n616) );
  INV_X1 U484 ( .A(KEYINPUT88), .ZN(n454) );
  NAND2_X1 U485 ( .A1(n379), .A2(n644), .ZN(n617) );
  XNOR2_X1 U486 ( .A(n380), .B(KEYINPUT107), .ZN(n379) );
  OR2_X1 U487 ( .A1(n554), .A2(n381), .ZN(n380) );
  XNOR2_X1 U488 ( .A(n584), .B(n420), .ZN(n596) );
  INV_X1 U489 ( .A(KEYINPUT76), .ZN(n420) );
  AND2_X1 U490 ( .A1(n662), .A2(n613), .ZN(n591) );
  XNOR2_X1 U491 ( .A(n537), .B(n724), .ZN(n705) );
  XNOR2_X1 U492 ( .A(n459), .B(n456), .ZN(n536) );
  XNOR2_X1 U493 ( .A(n495), .B(n487), .ZN(n403) );
  XNOR2_X1 U494 ( .A(n404), .B(n449), .ZN(n653) );
  NAND2_X1 U495 ( .A1(n652), .A2(KEYINPUT82), .ZN(n404) );
  XNOR2_X1 U496 ( .A(n455), .B(KEYINPUT40), .ZN(n737) );
  NAND2_X1 U497 ( .A1(n608), .A2(n644), .ZN(n455) );
  INV_X1 U498 ( .A(KEYINPUT35), .ZN(n438) );
  INV_X1 U499 ( .A(KEYINPUT32), .ZN(n385) );
  XNOR2_X1 U500 ( .A(n371), .B(KEYINPUT31), .ZN(n647) );
  AND2_X1 U501 ( .A1(n558), .A2(n542), .ZN(n646) );
  NOR2_X1 U502 ( .A1(n606), .A2(n593), .ZN(n642) );
  NOR2_X1 U503 ( .A1(n405), .A2(n383), .ZN(n382) );
  NAND2_X1 U504 ( .A1(n548), .A2(n384), .ZN(n383) );
  INV_X1 U505 ( .A(n549), .ZN(n384) );
  XNOR2_X1 U506 ( .A(n368), .B(KEYINPUT99), .ZN(n630) );
  AND2_X1 U507 ( .A1(n583), .A2(n548), .ZN(n369) );
  INV_X1 U508 ( .A(n658), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n466), .B(n359), .ZN(n465) );
  INV_X1 U510 ( .A(KEYINPUT126), .ZN(n414) );
  XNOR2_X1 U511 ( .A(n453), .B(n360), .ZN(n452) );
  AND2_X1 U512 ( .A1(n387), .A2(n554), .ZN(n351) );
  AND2_X1 U513 ( .A1(n364), .A2(n357), .ZN(n352) );
  XOR2_X1 U514 ( .A(G113), .B(G116), .Z(n353) );
  XNOR2_X1 U515 ( .A(KEYINPUT5), .B(KEYINPUT98), .ZN(n354) );
  OR2_X1 U516 ( .A1(n436), .A2(n429), .ZN(n355) );
  NAND2_X1 U517 ( .A1(n659), .A2(n603), .ZN(n356) );
  BUF_X1 U518 ( .A(n654), .Z(n405) );
  XNOR2_X1 U519 ( .A(n662), .B(KEYINPUT6), .ZN(n554) );
  INV_X1 U520 ( .A(G472), .ZN(n444) );
  INV_X1 U521 ( .A(n662), .ZN(n548) );
  AND2_X1 U522 ( .A1(n554), .A2(n450), .ZN(n357) );
  XOR2_X1 U523 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n358) );
  XOR2_X1 U524 ( .A(n627), .B(KEYINPUT110), .Z(n359) );
  XNOR2_X1 U525 ( .A(n373), .B(n390), .ZN(n725) );
  XNOR2_X1 U526 ( .A(n704), .B(KEYINPUT125), .ZN(n360) );
  NOR2_X1 U527 ( .A1(G952), .A2(n729), .ZN(n709) );
  INV_X1 U528 ( .A(n709), .ZN(n464) );
  INV_X1 U529 ( .A(KEYINPUT2), .ZN(n449) );
  XNOR2_X1 U530 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U531 ( .A1(n363), .A2(G478), .ZN(n453) );
  NAND2_X1 U532 ( .A1(n363), .A2(G472), .ZN(n466) );
  NAND2_X1 U533 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U534 ( .A(n655), .ZN(n361) );
  NOR2_X1 U535 ( .A1(n554), .A2(n361), .ZN(n362) );
  AND2_X2 U536 ( .A1(n349), .A2(n441), .ZN(n706) );
  BUF_X1 U537 ( .A(n386), .Z(n364) );
  XNOR2_X1 U538 ( .A(n366), .B(KEYINPUT22), .ZN(n386) );
  XNOR2_X1 U539 ( .A(n599), .B(n399), .ZN(n398) );
  NAND2_X1 U540 ( .A1(n706), .A2(G475), .ZN(n397) );
  NOR2_X2 U541 ( .A1(n556), .A2(n356), .ZN(n366) );
  NAND2_X1 U542 ( .A1(n351), .A2(n386), .ZN(n367) );
  NOR2_X1 U543 ( .A1(n647), .A2(n630), .ZN(n545) );
  INV_X1 U544 ( .A(n556), .ZN(n370) );
  NAND2_X1 U545 ( .A1(n370), .A2(n668), .ZN(n371) );
  XNOR2_X1 U546 ( .A(n372), .B(G122), .ZN(G24) );
  NAND2_X1 U547 ( .A1(n561), .A2(n372), .ZN(n562) );
  XNOR2_X2 U548 ( .A(n439), .B(n438), .ZN(n372) );
  XNOR2_X1 U549 ( .A(n373), .B(n530), .ZN(n413) );
  NAND2_X1 U550 ( .A1(n626), .A2(G472), .ZN(n374) );
  XNOR2_X1 U551 ( .A(n495), .B(n494), .ZN(n626) );
  XNOR2_X1 U552 ( .A(n611), .B(n610), .ZN(n377) );
  INV_X1 U553 ( .A(n613), .ZN(n381) );
  AND2_X1 U554 ( .A1(n364), .A2(n382), .ZN(n636) );
  NOR2_X1 U555 ( .A1(n617), .A2(n391), .ZN(n614) );
  XNOR2_X2 U556 ( .A(n392), .B(n491), .ZN(n504) );
  XNOR2_X2 U557 ( .A(n717), .B(KEYINPUT72), .ZN(n392) );
  XNOR2_X2 U558 ( .A(n482), .B(G107), .ZN(n717) );
  XNOR2_X1 U559 ( .A(n397), .B(n623), .ZN(n624) );
  INV_X1 U560 ( .A(n713), .ZN(n442) );
  AND2_X2 U561 ( .A1(n713), .A2(n449), .ZN(n443) );
  NAND2_X1 U562 ( .A1(n465), .A2(n464), .ZN(n463) );
  XNOR2_X1 U563 ( .A(n541), .B(n469), .ZN(n468) );
  XNOR2_X1 U564 ( .A(n406), .B(KEYINPUT53), .ZN(G75) );
  AND2_X1 U565 ( .A1(n691), .A2(n690), .ZN(n406) );
  NAND2_X1 U566 ( .A1(n600), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U567 ( .A1(n594), .A2(n642), .ZN(n600) );
  XNOR2_X1 U568 ( .A(n407), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X1 U569 ( .A(n415), .B(n414), .ZN(G63) );
  NAND2_X1 U570 ( .A1(n452), .A2(n464), .ZN(n415) );
  INV_X1 U571 ( .A(n649), .ZN(n421) );
  NOR2_X1 U572 ( .A1(n427), .A2(n426), .ZN(n425) );
  NOR2_X1 U573 ( .A1(n671), .A2(n430), .ZN(n426) );
  NOR2_X1 U574 ( .A1(n433), .A2(n429), .ZN(n427) );
  NAND2_X1 U575 ( .A1(n432), .A2(n436), .ZN(n431) );
  OR2_X1 U576 ( .A1(n626), .A2(n434), .ZN(n433) );
  NAND2_X1 U577 ( .A1(n440), .A2(n560), .ZN(n439) );
  XNOR2_X1 U578 ( .A(n557), .B(KEYINPUT34), .ZN(n440) );
  XNOR2_X2 U579 ( .A(n507), .B(n506), .ZN(n585) );
  XNOR2_X1 U580 ( .A(n503), .B(n716), .ZN(n446) );
  OR2_X1 U581 ( .A1(n713), .A2(n728), .ZN(n652) );
  XNOR2_X2 U582 ( .A(n574), .B(KEYINPUT45), .ZN(n713) );
  NOR2_X1 U583 ( .A1(n405), .A2(n451), .ZN(n450) );
  XNOR2_X1 U584 ( .A(n463), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U585 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U586 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U587 ( .A(n585), .ZN(n620) );
  XNOR2_X1 U588 ( .A(n350), .B(n692), .ZN(n694) );
  NOR2_X2 U589 ( .A1(n693), .A2(n622), .ZN(n507) );
  XNOR2_X1 U590 ( .A(n504), .B(n485), .ZN(n488) );
  AND2_X1 U591 ( .A1(G214), .A2(n492), .ZN(n470) );
  XNOR2_X1 U592 ( .A(KEYINPUT28), .B(n591), .ZN(n471) );
  OR2_X1 U593 ( .A1(n586), .A2(n644), .ZN(n594) );
  INV_X1 U594 ( .A(KEYINPUT25), .ZN(n539) );
  XNOR2_X1 U595 ( .A(n484), .B(KEYINPUT93), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U597 ( .A(n497), .B(n472), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U599 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n481) );
  XNOR2_X1 U600 ( .A(G143), .B(n486), .ZN(n473) );
  XNOR2_X1 U601 ( .A(n473), .B(G104), .ZN(n478) );
  XNOR2_X1 U602 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U603 ( .A(n533), .B(n479), .ZN(n521) );
  XNOR2_X1 U604 ( .A(n521), .B(KEYINPUT123), .ZN(n480) );
  XNOR2_X1 U605 ( .A(n481), .B(n480), .ZN(n623) );
  INV_X2 U606 ( .A(G953), .ZN(n729) );
  NAND2_X1 U607 ( .A1(G227), .A2(n729), .ZN(n483) );
  XNOR2_X1 U608 ( .A(n532), .B(n483), .ZN(n484) );
  XNOR2_X1 U609 ( .A(KEYINPUT71), .B(G469), .ZN(n489) );
  NAND2_X1 U610 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U611 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U612 ( .A(n517), .ZN(n622) );
  XNOR2_X1 U613 ( .A(n505), .B(KEYINPUT75), .ZN(n508) );
  NAND2_X1 U614 ( .A1(G210), .A2(n508), .ZN(n506) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n509) );
  NAND2_X1 U616 ( .A1(G234), .A2(G237), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n510), .B(KEYINPUT14), .ZN(n512) );
  NAND2_X1 U618 ( .A1(G952), .A2(n512), .ZN(n685) );
  NOR2_X1 U619 ( .A1(n685), .A2(G953), .ZN(n511) );
  XNOR2_X1 U620 ( .A(n511), .B(KEYINPUT90), .ZN(n578) );
  NAND2_X1 U621 ( .A1(n512), .A2(G902), .ZN(n513) );
  XNOR2_X1 U622 ( .A(KEYINPUT92), .B(n513), .ZN(n575) );
  XNOR2_X1 U623 ( .A(G898), .B(KEYINPUT91), .ZN(n712) );
  NAND2_X1 U624 ( .A1(G953), .A2(n712), .ZN(n720) );
  NOR2_X1 U625 ( .A1(n575), .A2(n720), .ZN(n514) );
  NOR2_X1 U626 ( .A1(n578), .A2(n514), .ZN(n515) );
  NAND2_X1 U627 ( .A1(G234), .A2(n517), .ZN(n518) );
  NAND2_X1 U628 ( .A1(n538), .A2(G221), .ZN(n520) );
  XNOR2_X1 U629 ( .A(KEYINPUT21), .B(n520), .ZN(n590) );
  INV_X1 U630 ( .A(n590), .ZN(n659) );
  NOR2_X1 U631 ( .A1(G902), .A2(n521), .ZN(n523) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(G475), .ZN(n522) );
  XNOR2_X1 U633 ( .A(n523), .B(n522), .ZN(n559) );
  XOR2_X1 U634 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n525) );
  XNOR2_X1 U635 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U636 ( .A1(G234), .A2(n729), .ZN(n529) );
  XOR2_X1 U637 ( .A(KEYINPUT8), .B(n529), .Z(n534) );
  NAND2_X1 U638 ( .A1(G217), .A2(n534), .ZN(n530) );
  NOR2_X1 U639 ( .A1(G902), .A2(n704), .ZN(n531) );
  XOR2_X1 U640 ( .A(G478), .B(n531), .Z(n558) );
  NOR2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n603) );
  XNOR2_X1 U642 ( .A(n533), .B(n532), .ZN(n724) );
  NAND2_X1 U643 ( .A1(G221), .A2(n534), .ZN(n535) );
  XNOR2_X1 U644 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U645 ( .A1(G217), .A2(n538), .ZN(n540) );
  INV_X1 U646 ( .A(n543), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n549), .B(KEYINPUT104), .ZN(n658) );
  XOR2_X1 U648 ( .A(KEYINPUT100), .B(n559), .Z(n542) );
  NOR2_X1 U649 ( .A1(n542), .A2(n558), .ZN(n644) );
  INV_X1 U650 ( .A(n594), .ZN(n676) );
  AND2_X1 U651 ( .A1(n592), .A2(n655), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n548), .A2(n553), .ZN(n668) );
  NOR2_X1 U653 ( .A1(n676), .A2(n545), .ZN(n546) );
  NOR2_X1 U654 ( .A1(n352), .A2(n546), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n547), .B(KEYINPUT105), .ZN(n551) );
  INV_X1 U656 ( .A(n567), .ZN(n552) );
  NOR2_X1 U657 ( .A1(n552), .A2(KEYINPUT66), .ZN(n550) );
  NOR2_X1 U658 ( .A1(n551), .A2(n550), .ZN(n564) );
  NAND2_X1 U659 ( .A1(n552), .A2(KEYINPUT66), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n556), .A2(n686), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n559), .A2(n558), .ZN(n595) );
  INV_X1 U662 ( .A(n595), .ZN(n560) );
  NAND2_X1 U663 ( .A1(n562), .A2(KEYINPUT44), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n564), .A2(n563), .ZN(n573) );
  INV_X1 U665 ( .A(KEYINPUT44), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n566), .A2(n567), .ZN(n569) );
  OR2_X1 U667 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n570) );
  NAND2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X2 U669 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U670 ( .A1(n729), .A2(n575), .ZN(n576) );
  NOR2_X1 U671 ( .A1(G900), .A2(n576), .ZN(n577) );
  NOR2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U673 ( .A(KEYINPUT81), .B(n579), .ZN(n588) );
  INV_X1 U674 ( .A(n588), .ZN(n580) );
  NOR2_X1 U675 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U676 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U677 ( .A(KEYINPUT38), .B(n620), .ZN(n672) );
  NAND2_X1 U678 ( .A1(n586), .A2(n608), .ZN(n587) );
  XNOR2_X1 U679 ( .A(n587), .B(KEYINPUT109), .ZN(n738) );
  NAND2_X1 U680 ( .A1(n543), .A2(n588), .ZN(n589) );
  NAND2_X1 U681 ( .A1(n471), .A2(n592), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n620), .A2(n595), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n641) );
  NAND2_X1 U684 ( .A1(n598), .A2(n641), .ZN(n599) );
  NOR2_X1 U685 ( .A1(KEYINPUT47), .A2(n600), .ZN(n601) );
  XNOR2_X1 U686 ( .A(n602), .B(KEYINPUT74), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n672), .A2(n671), .ZN(n675) );
  INV_X1 U688 ( .A(n603), .ZN(n674) );
  NOR2_X1 U689 ( .A1(n675), .A2(n674), .ZN(n605) );
  XNOR2_X1 U690 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n604) );
  XNOR2_X1 U691 ( .A(n605), .B(n604), .ZN(n687) );
  NOR2_X1 U692 ( .A1(n687), .A2(n606), .ZN(n607) );
  XOR2_X1 U693 ( .A(KEYINPUT42), .B(n607), .Z(n736) );
  NAND2_X1 U694 ( .A1(n736), .A2(n737), .ZN(n611) );
  XOR2_X1 U695 ( .A(KEYINPUT84), .B(KEYINPUT64), .Z(n609) );
  XOR2_X1 U696 ( .A(KEYINPUT36), .B(n614), .Z(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n649) );
  NOR2_X1 U698 ( .A1(n405), .A2(n617), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n618), .A2(n671), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT43), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n651) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT62), .ZN(n627) );
  XOR2_X1 U704 ( .A(G101), .B(n352), .Z(G3) );
  XOR2_X1 U705 ( .A(G104), .B(KEYINPUT111), .Z(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n644), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n629), .B(n628), .ZN(G6) );
  XOR2_X1 U708 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n632) );
  NAND2_X1 U709 ( .A1(n630), .A2(n646), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n632), .B(n631), .ZN(n633) );
  XOR2_X1 U711 ( .A(n633), .B(KEYINPUT112), .Z(n635) );
  XNOR2_X1 U712 ( .A(G107), .B(KEYINPUT26), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n635), .B(n634), .ZN(G9) );
  XOR2_X1 U714 ( .A(n636), .B(G110), .Z(G12) );
  XOR2_X1 U715 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n638) );
  NAND2_X1 U716 ( .A1(n642), .A2(n646), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U718 ( .A(G128), .B(n639), .ZN(G30) );
  XOR2_X1 U719 ( .A(G143), .B(KEYINPUT115), .Z(n640) );
  XNOR2_X1 U720 ( .A(n641), .B(n640), .ZN(G45) );
  NAND2_X1 U721 ( .A1(n642), .A2(n644), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(G146), .ZN(G48) );
  NAND2_X1 U723 ( .A1(n647), .A2(n644), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(G113), .ZN(G15) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n648), .B(G116), .ZN(G18) );
  XNOR2_X1 U727 ( .A(G125), .B(n649), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n650), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U729 ( .A(G140), .B(n651), .ZN(G42) );
  NOR2_X1 U730 ( .A1(G953), .A2(n653), .ZN(n691) );
  NOR2_X1 U731 ( .A1(n655), .A2(n405), .ZN(n657) );
  XNOR2_X1 U732 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n660), .Z(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(KEYINPUT117), .ZN(n664) );
  NOR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U739 ( .A(KEYINPUT119), .B(n666), .Z(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(n669), .Z(n670) );
  NOR2_X1 U742 ( .A1(n687), .A2(n670), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n686), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  XNOR2_X1 U750 ( .A(KEYINPUT120), .B(n683), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n706), .A2(G210), .ZN(n695) );
  XOR2_X1 U755 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n692) );
  XOR2_X1 U756 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n697) );
  XNOR2_X1 U757 ( .A(n698), .B(n697), .ZN(G51) );
  NAND2_X1 U758 ( .A1(n706), .A2(G469), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  NAND2_X1 U760 ( .A1(G217), .A2(n363), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n705), .B(n707), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n710) );
  XOR2_X1 U764 ( .A(KEYINPUT61), .B(n710), .Z(n711) );
  NOR2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U766 ( .A1(G953), .A2(n713), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n723) );
  XOR2_X1 U768 ( .A(KEYINPUT127), .B(n716), .Z(n719) );
  XNOR2_X1 U769 ( .A(n717), .B(G101), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U772 ( .A(n723), .B(n722), .ZN(G69) );
  XOR2_X1 U773 ( .A(n725), .B(n724), .Z(n726) );
  XNOR2_X1 U774 ( .A(n727), .B(n726), .ZN(n731) );
  XNOR2_X1 U775 ( .A(n731), .B(n728), .ZN(n730) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n735) );
  XNOR2_X1 U777 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U778 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U779 ( .A1(G953), .A2(n733), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n735), .A2(n734), .ZN(G72) );
  XOR2_X1 U781 ( .A(n365), .B(G119), .Z(G21) );
  XNOR2_X1 U782 ( .A(G137), .B(n736), .ZN(G39) );
  XNOR2_X1 U783 ( .A(G131), .B(n737), .ZN(G33) );
  XOR2_X1 U784 ( .A(G134), .B(n738), .Z(n739) );
  XNOR2_X1 U785 ( .A(KEYINPUT116), .B(n739), .ZN(G36) );
endmodule

