

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U555 ( .A(n609), .B(KEYINPUT31), .ZN(n668) );
  OR2_X2 U556 ( .A1(n608), .A2(n607), .ZN(n609) );
  OR2_X1 U557 ( .A1(n602), .A2(n601), .ZN(n603) );
  BUF_X1 U558 ( .A(n899), .Z(n522) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(n523), .Z(n899) );
  XNOR2_X1 U560 ( .A(n682), .B(KEYINPUT104), .ZN(n683) );
  NOR2_X1 U561 ( .A1(n697), .A2(n696), .ZN(n698) );
  AND2_X1 U562 ( .A1(n683), .A2(n705), .ZN(n687) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G651), .A2(n588), .ZN(n803) );
  AND2_X1 U565 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U566 ( .A1(n534), .A2(n533), .ZN(G160) );
  NAND2_X1 U567 ( .A1(n522), .A2(G137), .ZN(n524) );
  XNOR2_X1 U568 ( .A(n524), .B(KEYINPUT66), .ZN(n526) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U570 ( .A1(G113), .A2(n894), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U572 ( .A(n527), .B(KEYINPUT67), .ZN(n534) );
  XOR2_X1 U573 ( .A(KEYINPUT65), .B(KEYINPUT23), .Z(n529) );
  INV_X1 U574 ( .A(G2105), .ZN(n530) );
  AND2_X1 U575 ( .A1(n530), .A2(G2104), .ZN(n897) );
  NAND2_X1 U576 ( .A1(G101), .A2(n897), .ZN(n528) );
  XOR2_X1 U577 ( .A(n529), .B(n528), .Z(n532) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n530), .ZN(n893) );
  NAND2_X1 U579 ( .A1(G125), .A2(n893), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G138), .A2(n522), .ZN(n536) );
  NAND2_X1 U581 ( .A1(G102), .A2(n897), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U583 ( .A(n537), .B(KEYINPUT92), .ZN(n541) );
  NAND2_X1 U584 ( .A1(G126), .A2(n893), .ZN(n539) );
  NAND2_X1 U585 ( .A1(G114), .A2(n894), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U587 ( .A1(n541), .A2(n540), .ZN(G164) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n808) );
  NAND2_X1 U589 ( .A1(n808), .A2(G89), .ZN(n542) );
  XNOR2_X1 U590 ( .A(n542), .B(KEYINPUT4), .ZN(n545) );
  INV_X1 U591 ( .A(G651), .ZN(n547) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n588) );
  OR2_X1 U593 ( .A1(n547), .A2(n588), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n543), .Z(n805) );
  NAND2_X1 U595 ( .A1(G76), .A2(n805), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U597 ( .A(n546), .B(KEYINPUT5), .ZN(n553) );
  NOR2_X1 U598 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n548), .Z(n809) );
  NAND2_X1 U600 ( .A1(G63), .A2(n809), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G51), .A2(n803), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U604 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U605 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U606 ( .A1(G64), .A2(n809), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G52), .A2(n803), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U609 ( .A1(G77), .A2(n805), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n808), .A2(G90), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U613 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U614 ( .A1(n803), .A2(G53), .ZN(n568) );
  NAND2_X1 U615 ( .A1(n809), .A2(G65), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G78), .A2(n805), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U618 ( .A1(n808), .A2(G91), .ZN(n564) );
  XOR2_X1 U619 ( .A(KEYINPUT70), .B(n564), .Z(n565) );
  NOR2_X1 U620 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U622 ( .A(KEYINPUT71), .B(n569), .Z(G299) );
  NAND2_X1 U623 ( .A1(G88), .A2(n808), .ZN(n571) );
  NAND2_X1 U624 ( .A1(G75), .A2(n805), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U626 ( .A1(G62), .A2(n809), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G50), .A2(n803), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U629 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U630 ( .A(KEYINPUT82), .B(n576), .Z(G303) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(n805), .A2(G73), .ZN(n577) );
  XNOR2_X1 U633 ( .A(n577), .B(KEYINPUT2), .ZN(n584) );
  NAND2_X1 U634 ( .A1(G86), .A2(n808), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G61), .A2(n809), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G48), .A2(n803), .ZN(n580) );
  XNOR2_X1 U638 ( .A(KEYINPUT81), .B(n580), .ZN(n581) );
  NOR2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U641 ( .A1(G49), .A2(n803), .ZN(n586) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U644 ( .A1(n809), .A2(n587), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n588), .A2(G87), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G85), .A2(n808), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G72), .A2(n805), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U650 ( .A1(G60), .A2(n809), .ZN(n593) );
  XNOR2_X1 U651 ( .A(KEYINPUT69), .B(n593), .ZN(n594) );
  NOR2_X1 U652 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U653 ( .A1(n803), .A2(G47), .ZN(n596) );
  NAND2_X1 U654 ( .A1(n597), .A2(n596), .ZN(G290) );
  NOR2_X1 U655 ( .A1(G1384), .A2(G164), .ZN(n598) );
  XOR2_X1 U656 ( .A(n598), .B(KEYINPUT64), .Z(n727) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n729) );
  NOR2_X2 U658 ( .A1(n727), .A2(n729), .ZN(n637) );
  INV_X1 U659 ( .A(n637), .ZN(n622) );
  NOR2_X1 U660 ( .A1(G2084), .A2(n622), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G8), .A2(n599), .ZN(n663) );
  NAND2_X1 U662 ( .A1(n622), .A2(G8), .ZN(n705) );
  NOR2_X1 U663 ( .A1(G1966), .A2(n705), .ZN(n602) );
  INV_X1 U664 ( .A(n599), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G8), .A2(n600), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n603), .B(KEYINPUT30), .ZN(n604) );
  NOR2_X1 U667 ( .A1(G168), .A2(n604), .ZN(n608) );
  INV_X1 U668 ( .A(G1961), .ZN(n962) );
  NAND2_X1 U669 ( .A1(n622), .A2(n962), .ZN(n606) );
  XNOR2_X1 U670 ( .A(G2078), .B(KEYINPUT25), .ZN(n931) );
  NAND2_X1 U671 ( .A1(n637), .A2(n931), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n606), .A2(n605), .ZN(n658) );
  NOR2_X1 U673 ( .A1(G171), .A2(n658), .ZN(n607) );
  INV_X1 U674 ( .A(G299), .ZN(n815) );
  NAND2_X1 U675 ( .A1(n637), .A2(G2072), .ZN(n610) );
  XNOR2_X1 U676 ( .A(n610), .B(KEYINPUT27), .ZN(n612) );
  INV_X1 U677 ( .A(G1956), .ZN(n950) );
  NOR2_X1 U678 ( .A1(n950), .A2(n637), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n653) );
  NAND2_X1 U680 ( .A1(n815), .A2(n653), .ZN(n651) );
  NAND2_X1 U681 ( .A1(G66), .A2(n809), .ZN(n619) );
  NAND2_X1 U682 ( .A1(G92), .A2(n808), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G79), .A2(n805), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G54), .A2(n803), .ZN(n615) );
  XNOR2_X1 U686 ( .A(KEYINPUT75), .B(n615), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT15), .ZN(n915) );
  NAND2_X1 U690 ( .A1(G2067), .A2(n637), .ZN(n621) );
  XOR2_X1 U691 ( .A(KEYINPUT98), .B(n621), .Z(n624) );
  AND2_X1 U692 ( .A1(n622), .A2(G1348), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U694 ( .A1(n915), .A2(n625), .ZN(n649) );
  NAND2_X1 U695 ( .A1(n915), .A2(n625), .ZN(n647) );
  NAND2_X1 U696 ( .A1(G81), .A2(n808), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT12), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT74), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G68), .A2(n805), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT13), .B(n630), .Z(n634) );
  NAND2_X1 U702 ( .A1(G56), .A2(n809), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT14), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT73), .ZN(n633) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n803), .A2(G43), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n1019) );
  AND2_X1 U708 ( .A1(n637), .A2(G1996), .ZN(n639) );
  INV_X1 U709 ( .A(KEYINPUT26), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n642) );
  INV_X1 U711 ( .A(n639), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n640), .A2(KEYINPUT26), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n622), .A2(G1341), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  OR2_X1 U716 ( .A1(n1019), .A2(n645), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n652), .B(KEYINPUT99), .ZN(n656) );
  OR2_X1 U721 ( .A1(n815), .A2(n653), .ZN(n654) );
  XOR2_X1 U722 ( .A(KEYINPUT28), .B(n654), .Z(n655) );
  NOR2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT29), .B(n657), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n658), .A2(G171), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n670) );
  AND2_X1 U727 ( .A1(n668), .A2(n670), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n602), .A2(n661), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n688) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n705), .ZN(n665) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n622), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U733 ( .A1(G303), .A2(n666), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT100), .ZN(n671) );
  AND2_X1 U735 ( .A1(n668), .A2(n671), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n674) );
  INV_X1 U737 ( .A(n671), .ZN(n672) );
  OR2_X1 U738 ( .A1(n672), .A2(G286), .ZN(n673) );
  AND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U740 ( .A1(G8), .A2(n675), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n676) );
  XNOR2_X1 U742 ( .A(n677), .B(n676), .ZN(n690) );
  NAND2_X1 U743 ( .A1(n688), .A2(n690), .ZN(n681) );
  NOR2_X1 U744 ( .A1(G303), .A2(G2090), .ZN(n678) );
  XOR2_X1 U745 ( .A(KEYINPUT103), .B(n678), .Z(n679) );
  NAND2_X1 U746 ( .A1(G8), .A2(n679), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  INV_X1 U748 ( .A(n705), .ZN(n695) );
  NOR2_X1 U749 ( .A1(G1981), .A2(G305), .ZN(n684) );
  XOR2_X1 U750 ( .A(n684), .B(KEYINPUT24), .Z(n685) );
  NOR2_X1 U751 ( .A1(n705), .A2(n685), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n710) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  AND2_X1 U754 ( .A1(n688), .A2(n1005), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n694) );
  INV_X1 U756 ( .A(n1005), .ZN(n692) );
  NOR2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n700) );
  NOR2_X1 U758 ( .A1(G303), .A2(G1971), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n700), .A2(n691), .ZN(n1006) );
  OR2_X1 U760 ( .A1(n692), .A2(n1006), .ZN(n693) );
  AND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n695), .A2(KEYINPUT102), .ZN(n696) );
  NOR2_X1 U763 ( .A1(KEYINPUT33), .A2(n698), .ZN(n707) );
  INV_X1 U764 ( .A(KEYINPUT102), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n699), .A2(n700), .ZN(n703) );
  NAND2_X1 U766 ( .A1(n700), .A2(KEYINPUT33), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n701), .A2(KEYINPUT102), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U771 ( .A(G1981), .B(G305), .Z(n1015) );
  NAND2_X1 U772 ( .A1(n708), .A2(n1015), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n745) );
  NAND2_X1 U774 ( .A1(G131), .A2(n522), .ZN(n712) );
  NAND2_X1 U775 ( .A1(G95), .A2(n897), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U777 ( .A1(G119), .A2(n893), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G107), .A2(n894), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n879) );
  XOR2_X1 U781 ( .A(KEYINPUT96), .B(G1991), .Z(n933) );
  NOR2_X1 U782 ( .A1(n879), .A2(n933), .ZN(n717) );
  XOR2_X1 U783 ( .A(KEYINPUT97), .B(n717), .Z(n726) );
  INV_X1 U784 ( .A(G1996), .ZN(n928) );
  NAND2_X1 U785 ( .A1(G105), .A2(n897), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n718), .B(KEYINPUT38), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n522), .A2(G141), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U789 ( .A1(G129), .A2(n893), .ZN(n722) );
  NAND2_X1 U790 ( .A1(G117), .A2(n894), .ZN(n721) );
  NAND2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n906) );
  NOR2_X1 U793 ( .A1(n928), .A2(n906), .ZN(n725) );
  NOR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n748) );
  XOR2_X1 U795 ( .A(G1986), .B(G290), .Z(n1009) );
  NAND2_X1 U796 ( .A1(n748), .A2(n1009), .ZN(n730) );
  INV_X1 U797 ( .A(n727), .ZN(n728) );
  NOR2_X1 U798 ( .A1(n729), .A2(n728), .ZN(n755) );
  NAND2_X1 U799 ( .A1(n730), .A2(n755), .ZN(n743) );
  XNOR2_X1 U800 ( .A(KEYINPUT36), .B(KEYINPUT95), .ZN(n742) );
  NAND2_X1 U801 ( .A1(G140), .A2(n522), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G104), .A2(n897), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U804 ( .A(KEYINPUT34), .B(n733), .ZN(n739) );
  NAND2_X1 U805 ( .A1(n893), .A2(G128), .ZN(n734) );
  XOR2_X1 U806 ( .A(KEYINPUT93), .B(n734), .Z(n736) );
  NAND2_X1 U807 ( .A1(n894), .A2(G116), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U809 ( .A(n737), .B(KEYINPUT35), .Z(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U811 ( .A(KEYINPUT94), .B(n740), .Z(n741) );
  XOR2_X1 U812 ( .A(n742), .B(n741), .Z(n910) );
  XOR2_X1 U813 ( .A(KEYINPUT37), .B(G2067), .Z(n746) );
  AND2_X1 U814 ( .A1(n910), .A2(n746), .ZN(n987) );
  NAND2_X1 U815 ( .A1(n987), .A2(n755), .ZN(n747) );
  AND2_X1 U816 ( .A1(n743), .A2(n747), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n762) );
  NOR2_X1 U818 ( .A1(n746), .A2(n910), .ZN(n995) );
  NAND2_X1 U819 ( .A1(n995), .A2(n755), .ZN(n760) );
  INV_X1 U820 ( .A(n747), .ZN(n758) );
  AND2_X1 U821 ( .A1(n928), .A2(n906), .ZN(n979) );
  INV_X1 U822 ( .A(n748), .ZN(n991) );
  NAND2_X1 U823 ( .A1(n933), .A2(n879), .ZN(n749) );
  XOR2_X1 U824 ( .A(KEYINPUT106), .B(n749), .Z(n982) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n750) );
  XOR2_X1 U826 ( .A(n750), .B(KEYINPUT105), .Z(n751) );
  NOR2_X1 U827 ( .A1(n982), .A2(n751), .ZN(n752) );
  NOR2_X1 U828 ( .A1(n991), .A2(n752), .ZN(n753) );
  NOR2_X1 U829 ( .A1(n979), .A2(n753), .ZN(n754) );
  XNOR2_X1 U830 ( .A(KEYINPUT39), .B(n754), .ZN(n756) );
  NAND2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n757) );
  OR2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U833 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U835 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U836 ( .A(G2451), .B(G2443), .ZN(n773) );
  XOR2_X1 U837 ( .A(G2446), .B(G2430), .Z(n765) );
  XNOR2_X1 U838 ( .A(KEYINPUT108), .B(G2438), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n765), .B(n764), .ZN(n769) );
  XOR2_X1 U840 ( .A(G2435), .B(G2454), .Z(n767) );
  XNOR2_X1 U841 ( .A(G1348), .B(G1341), .ZN(n766) );
  XNOR2_X1 U842 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U843 ( .A(n769), .B(n768), .Z(n771) );
  XNOR2_X1 U844 ( .A(KEYINPUT107), .B(G2427), .ZN(n770) );
  XNOR2_X1 U845 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U846 ( .A(n773), .B(n772), .ZN(n774) );
  AND2_X1 U847 ( .A1(n774), .A2(G14), .ZN(G401) );
  AND2_X1 U848 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  INV_X1 U851 ( .A(G57), .ZN(G237) );
  INV_X1 U852 ( .A(G108), .ZN(G238) );
  INV_X1 U853 ( .A(G120), .ZN(G236) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U855 ( .A(n775), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U856 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n777) );
  INV_X1 U857 ( .A(G223), .ZN(n848) );
  NAND2_X1 U858 ( .A1(G567), .A2(n848), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n777), .B(n776), .ZN(G234) );
  INV_X1 U860 ( .A(G860), .ZN(n802) );
  OR2_X1 U861 ( .A1(n1019), .A2(n802), .ZN(G153) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  INV_X1 U863 ( .A(n915), .ZN(n1018) );
  INV_X1 U864 ( .A(G868), .ZN(n785) );
  NAND2_X1 U865 ( .A1(n1018), .A2(n785), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT76), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G868), .A2(G301), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(G284) );
  NAND2_X1 U869 ( .A1(G286), .A2(G868), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G299), .A2(n785), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U872 ( .A1(n802), .A2(G559), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n783), .A2(n915), .ZN(n784) );
  XNOR2_X1 U874 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U875 ( .A1(G559), .A2(n785), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n915), .A2(n786), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(KEYINPUT77), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n1019), .A2(G868), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U880 ( .A1(G123), .A2(n893), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT18), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G99), .A2(n897), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT79), .B(n791), .Z(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G135), .A2(n522), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n794), .B(KEYINPUT78), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n894), .A2(G111), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n983) );
  XNOR2_X1 U890 ( .A(n983), .B(G2096), .ZN(n800) );
  INV_X1 U891 ( .A(G2100), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(G156) );
  NAND2_X1 U893 ( .A1(G559), .A2(n915), .ZN(n801) );
  XOR2_X1 U894 ( .A(n1019), .B(n801), .Z(n824) );
  NAND2_X1 U895 ( .A1(n802), .A2(n824), .ZN(n814) );
  NAND2_X1 U896 ( .A1(G55), .A2(n803), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n804), .B(KEYINPUT80), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G80), .A2(n805), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G93), .A2(n808), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G67), .A2(n809), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n826) );
  XOR2_X1 U904 ( .A(n814), .B(n826), .Z(G145) );
  INV_X1 U905 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U906 ( .A(n815), .B(G166), .ZN(n823) );
  XOR2_X1 U907 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n816) );
  XNOR2_X1 U908 ( .A(G288), .B(n816), .ZN(n817) );
  XNOR2_X1 U909 ( .A(KEYINPUT85), .B(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(G305), .B(KEYINPUT84), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n826), .B(n820), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(G290), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n823), .B(n822), .ZN(n914) );
  XNOR2_X1 U915 ( .A(n824), .B(n914), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n825), .A2(G868), .ZN(n828) );
  OR2_X1 U917 ( .A1(G868), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(G295) );
  NAND2_X1 U919 ( .A1(G2078), .A2(G2084), .ZN(n830) );
  XOR2_X1 U920 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n829) );
  XNOR2_X1 U921 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G2090), .A2(n831), .ZN(n832) );
  XNOR2_X1 U923 ( .A(KEYINPUT21), .B(n832), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n833), .A2(G2072), .ZN(n834) );
  XOR2_X1 U925 ( .A(KEYINPUT87), .B(n834), .Z(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U927 ( .A1(G236), .A2(G238), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G69), .A2(n835), .ZN(n836) );
  NOR2_X1 U929 ( .A1(n836), .A2(G237), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(KEYINPUT89), .ZN(n852) );
  NAND2_X1 U931 ( .A1(G567), .A2(n852), .ZN(n843) );
  NOR2_X1 U932 ( .A1(G220), .A2(G219), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT22), .B(n838), .Z(n839) );
  NOR2_X1 U934 ( .A1(G218), .A2(n839), .ZN(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT88), .B(n840), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n841), .A2(G96), .ZN(n853) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n853), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT90), .B(n844), .Z(G319) );
  INV_X1 U940 ( .A(G319), .ZN(n846) );
  NAND2_X1 U941 ( .A1(G661), .A2(G483), .ZN(n845) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U943 ( .A(KEYINPUT91), .B(n847), .Z(n851) );
  NAND2_X1 U944 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n848), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U947 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(G188) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1976), .B(G1981), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1966), .B(G1956), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(n864), .B(G2474), .Z(n866) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT41), .B(G1986), .Z(n868) );
  XNOR2_X1 U970 ( .A(G1961), .B(G1971), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n893), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G136), .A2(n522), .ZN(n872) );
  XOR2_X1 U976 ( .A(KEYINPUT109), .B(n872), .Z(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G112), .A2(n894), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G100), .A2(n897), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(G162) );
  XOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n881) );
  XNOR2_X1 U983 ( .A(n879), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U985 ( .A(n882), .B(n983), .Z(n892) );
  NAND2_X1 U986 ( .A1(G139), .A2(n522), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G103), .A2(n897), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n885), .Z(n890) );
  NAND2_X1 U990 ( .A1(G127), .A2(n893), .ZN(n887) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n886) );
  NAND2_X1 U992 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n997) );
  XNOR2_X1 U995 ( .A(G164), .B(n997), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n892), .B(n891), .ZN(n909) );
  NAND2_X1 U997 ( .A1(G130), .A2(n893), .ZN(n896) );
  NAND2_X1 U998 ( .A1(G118), .A2(n894), .ZN(n895) );
  NAND2_X1 U999 ( .A1(n896), .A2(n895), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n897), .A2(G106), .ZN(n898) );
  XNOR2_X1 U1001 ( .A(n898), .B(KEYINPUT110), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n522), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1004 ( .A(KEYINPUT45), .B(n902), .Z(n903) );
  NOR2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(G162), .B(n905), .ZN(n907) );
  XOR2_X1 U1007 ( .A(n907), .B(n906), .Z(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(G160), .B(n910), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n913), .ZN(G395) );
  XOR2_X1 U1012 ( .A(KEYINPUT113), .B(n914), .Z(n917) );
  XNOR2_X1 U1013 ( .A(n915), .B(G286), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n1019), .B(G171), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n920), .ZN(G397) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n923), .ZN(n924) );
  AND2_X1 U1022 ( .A1(n924), .A2(G319), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1027 ( .A(G2084), .B(G34), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT54), .ZN(n946) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n943) );
  XOR2_X1 U1030 ( .A(G2072), .B(G33), .Z(n930) );
  XNOR2_X1 U1031 ( .A(n928), .B(G32), .ZN(n929) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G27), .B(n931), .ZN(n938) );
  XOR2_X1 U1034 ( .A(G2067), .B(G26), .Z(n932) );
  NAND2_X1 U1035 ( .A1(n932), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT119), .B(n933), .ZN(n934) );
  XNOR2_X1 U1037 ( .A(G25), .B(n934), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1043 ( .A(KEYINPUT120), .B(n944), .Z(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1045 ( .A(KEYINPUT121), .B(n947), .Z(n948) );
  NOR2_X1 U1046 ( .A1(G29), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT55), .B(n949), .ZN(n1034) );
  XNOR2_X1 U1048 ( .A(G20), .B(n950), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1053 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1054 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1056 ( .A(KEYINPUT60), .B(n958), .Z(n960) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G21), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(KEYINPUT124), .B(n961), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n962), .B(G5), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G1971), .B(G22), .Z(n965) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1066 ( .A(KEYINPUT126), .B(n968), .Z(n970) );
  XNOR2_X1 U1067 ( .A(G1986), .B(G24), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1069 ( .A(KEYINPUT58), .B(n971), .Z(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n974), .B(KEYINPUT61), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT123), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n977), .ZN(n1032) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT51), .B(n980), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(n981), .B(KEYINPUT117), .ZN(n993) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1080 ( .A(KEYINPUT115), .B(n984), .Z(n986) );
  XNOR2_X1 U1081 ( .A(G160), .B(G2084), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1084 ( .A(KEYINPUT116), .B(n989), .Z(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT118), .B(n996), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(G2072), .B(n997), .Z(n999) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(n1003), .B(KEYINPUT52), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(G29), .ZN(n1030) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  AND2_X1 U1097 ( .A1(G303), .A2(G1971), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G171), .B(G1961), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G1956), .B(G299), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1025) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G168), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT57), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1018), .B(G1348), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1019), .B(G1341), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT122), .B(n1026), .Z(n1028) );
  XNOR2_X1 U1113 ( .A(G16), .B(KEYINPUT56), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(n1035), .B(KEYINPUT127), .ZN(n1036) );
  XNOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1036), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

