//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT39), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT77), .B1(new_n208), .B2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(G141gat), .B2(new_n210), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n208), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n203), .B(new_n206), .C1(new_n214), .C2(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G127gat), .B(G134gat), .Z(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n222));
  INV_X1    g021(.A(G113gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G120gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n226));
  AOI211_X1 g025(.A(KEYINPUT1), .B(new_n219), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n224), .B2(new_n221), .ZN(new_n229));
  INV_X1    g028(.A(G127gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n229), .B(new_n231), .C1(KEYINPUT68), .C2(new_n219), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n232), .B(new_n233), .ZN(new_n239));
  INV_X1    g038(.A(new_n227), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(new_n216), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT81), .B(new_n238), .C1(new_n242), .C2(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n216), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n216), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n252));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT78), .Z(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n202), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT88), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n236), .A2(new_n247), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n242), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n254), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n202), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT87), .Z(new_n270));
  NAND3_X1  g069(.A1(new_n257), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT40), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT74), .B(G218gat), .Z(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n274), .B1(new_n277), .B2(KEYINPUT22), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT27), .B(G183gat), .Z(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n287), .A2(new_n288), .A3(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n287), .B2(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT65), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n281), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n296), .B(new_n297), .C1(G183gat), .C2(G190gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT64), .B(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT23), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n294), .A2(new_n298), .A3(new_n283), .A4(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n292), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n283), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  NOR4_X1   g107(.A1(new_n305), .A2(new_n307), .A3(new_n303), .A4(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n281), .B1(new_n310), .B2(KEYINPUT24), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n312));
  OAI221_X1 g111(.A(new_n297), .B1(G183gat), .B2(G190gat), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n294), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n291), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n315), .B2(KEYINPUT29), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n318), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n280), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n280), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT76), .B(new_n316), .C1(new_n315), .C2(KEYINPUT29), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n317), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n323), .A2(new_n328), .A3(new_n332), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT30), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n323), .A2(new_n337), .A3(new_n328), .A4(new_n332), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n257), .A2(new_n265), .A3(KEYINPUT40), .A4(new_n270), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n248), .A2(new_n237), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n254), .B1(new_n241), .B2(new_n245), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n218), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n254), .B1(new_n242), .B2(new_n261), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n241), .A2(new_n216), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n263), .B1(new_n349), .B2(new_n248), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n345), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n243), .A3(new_n250), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT89), .B1(new_n358), .B2(new_n270), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n360));
  INV_X1    g159(.A(new_n270), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n360), .B(new_n361), .C1(new_n353), .C2(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n273), .A2(new_n339), .A3(new_n340), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n336), .A2(new_n338), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n359), .B2(new_n362), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(KEYINPUT90), .A3(new_n340), .A4(new_n273), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT31), .B(G50gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G22gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n373), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT29), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n326), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n244), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n247), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n384), .A2(new_n218), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n380), .B1(new_n388), .B2(KEYINPUT84), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n384), .A2(KEYINPUT84), .A3(new_n218), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n389), .A2(new_n390), .B1(G228gat), .B2(G233gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n377), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n381), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n385), .B(KEYINPUT85), .ZN(new_n395));
  INV_X1    g194(.A(new_n377), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n333), .B1(new_n329), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(KEYINPUT37), .B2(new_n329), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n322), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n280), .B1(new_n405), .B2(new_n319), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n325), .A2(new_n317), .A3(new_n327), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT37), .B1(new_n407), .B2(new_n326), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n335), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n269), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT6), .B(new_n412), .C1(new_n353), .C2(new_n357), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT94), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT80), .B1(new_n346), .B2(KEYINPUT5), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n350), .A2(new_n348), .A3(new_n351), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n344), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n356), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT6), .A4(new_n412), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT6), .B1(new_n358), .B2(new_n269), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT91), .B1(new_n363), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n360), .B1(new_n421), .B2(new_n361), .ZN(new_n429));
  INV_X1    g228(.A(new_n362), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT91), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n411), .B(new_n426), .C1(new_n428), .C2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n370), .A2(new_n398), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n241), .A2(new_n315), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n241), .A2(new_n315), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT34), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n436), .A2(new_n437), .B1(G227gat), .B2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n443), .A2(KEYINPUT72), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n435), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n436), .A2(G227gat), .A3(G233gat), .A4(new_n437), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(KEYINPUT32), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n450), .A2(KEYINPUT32), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n449), .A2(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(KEYINPUT71), .A3(new_n453), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n446), .A2(new_n456), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT34), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n444), .B1(new_n443), .B2(KEYINPUT72), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT73), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n467), .A2(new_n435), .B1(new_n457), .B2(new_n458), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n464), .A3(new_n456), .A4(new_n460), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(KEYINPUT36), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n414), .A2(new_n415), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n421), .A2(new_n475), .A3(new_n412), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n412), .B1(new_n353), .B2(new_n357), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n427), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n339), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n470), .B(new_n473), .C1(new_n480), .C2(new_n398), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n434), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n424), .B1(new_n417), .B2(new_n423), .ZN(new_n484));
  INV_X1    g283(.A(new_n425), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n432), .A2(new_n428), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  AND4_X1   g286(.A1(new_n487), .A2(new_n471), .A3(new_n367), .A4(new_n398), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n423), .A3(new_n417), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(new_n367), .A3(new_n398), .A4(new_n471), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n486), .A2(new_n488), .B1(new_n490), .B2(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT14), .B(G29gat), .Z(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G43gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(G43gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n504), .B2(new_n499), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT95), .B(KEYINPUT15), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n508), .A2(new_n497), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n493), .B(new_n503), .C1(new_n509), .C2(new_n502), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(G8gat), .Z(new_n515));
  AOI21_X1  g314(.A(new_n502), .B1(new_n508), .B2(new_n497), .ZN(new_n516));
  INV_X1    g315(.A(new_n503), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT17), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n510), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n515), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT18), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n522), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n523), .B(KEYINPUT13), .Z(new_n530));
  AOI22_X1  g329(.A1(new_n524), .A2(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n519), .A2(new_n523), .A3(new_n522), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G197gat), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT11), .B(G169gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT12), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(KEYINPUT98), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n532), .A2(new_n543), .A3(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n540), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n526), .A3(new_n531), .A4(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n483), .A2(new_n492), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT41), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  NOR2_X1   g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(KEYINPUT8), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(new_n552), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n550), .B1(new_n527), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n510), .A2(new_n518), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(KEYINPUT102), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT103), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(KEYINPUT103), .A3(new_n564), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G190gat), .B(G218gat), .Z(new_n570));
  OR2_X1    g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G134gat), .B(G162gat), .Z(new_n572));
  NOR2_X1   g371(.A1(new_n549), .A2(KEYINPUT41), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT104), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n569), .B2(new_n570), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(KEYINPUT104), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT105), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(new_n577), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g384(.A(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G57gat), .ZN(new_n587));
  INV_X1    g386(.A(G57gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT99), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n585), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT100), .B(G57gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n587), .B1(new_n600), .B2(new_n586), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n585), .A2(G71gat), .A3(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT21), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G127gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n599), .A2(new_n609), .A3(new_n604), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n599), .B2(new_n604), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n520), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n608), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n618), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n584), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n588), .A2(G64gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n586), .A2(G57gat), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT9), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n596), .B1(new_n630), .B2(new_n595), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n604), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n561), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n599), .A2(new_n558), .A3(new_n604), .A4(new_n560), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(KEYINPUT101), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n599), .A2(new_n609), .A3(new_n604), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT106), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT107), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647));
  AOI211_X1 g446(.A(new_n647), .B(new_n644), .C1(new_n637), .C2(new_n641), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n634), .B2(new_n636), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n627), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n650), .B(new_n627), .C1(new_n642), .C2(new_n645), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n623), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n548), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n489), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n339), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n548), .A2(new_n655), .ZN(new_n662));
  OAI21_X1  g461(.A(G8gat), .B1(new_n662), .B2(new_n367), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  MUX2_X1   g463(.A(new_n661), .B(new_n664), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g464(.A1(new_n473), .A2(new_n470), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT108), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n471), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n662), .B2(new_n670), .ZN(G1326gat));
  INV_X1    g470(.A(new_n398), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n656), .A2(KEYINPUT109), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n662), .B2(new_n398), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n547), .A2(new_n541), .ZN(new_n680));
  INV_X1    g479(.A(new_n654), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n584), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT91), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n687), .A2(new_n431), .B1(new_n416), .B2(new_n425), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n672), .B1(new_n688), .B2(new_n411), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n481), .B1(new_n689), .B2(new_n370), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n680), .B(new_n684), .C1(new_n690), .C2(new_n491), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(G29gat), .A3(new_n489), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT45), .Z(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n491), .B1(new_n434), .B2(new_n482), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n683), .ZN(new_n696));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n584), .C1(new_n690), .C2(new_n491), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n680), .A2(KEYINPUT110), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n547), .B2(new_n541), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n682), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n698), .A2(new_n657), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n693), .B1(new_n494), .B2(new_n705), .ZN(G1328gat));
  NOR3_X1   g505(.A1(new_n691), .A2(G36gat), .A3(new_n367), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n698), .A2(new_n339), .A3(new_n704), .ZN(new_n709));
  INV_X1    g508(.A(G36gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(G1329gat));
  NOR2_X1   g510(.A1(new_n669), .A2(G43gat), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n548), .A2(KEYINPUT111), .A3(new_n684), .A4(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  INV_X1    g513(.A(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n691), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n713), .A2(new_n716), .B1(KEYINPUT112), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n666), .A3(new_n697), .A4(new_n704), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(KEYINPUT47), .A3(G43gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n713), .A2(new_n716), .ZN(new_n722));
  INV_X1    g521(.A(new_n667), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n696), .A2(new_n723), .A3(new_n697), .A4(new_n704), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n722), .A2(KEYINPUT112), .B1(G43gat), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n725), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g525(.A1(new_n398), .A2(new_n498), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n704), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n498), .B1(new_n691), .B2(new_n398), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n728), .B2(new_n729), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  NOR4_X1   g532(.A1(new_n695), .A2(new_n623), .A3(new_n681), .A4(new_n702), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n657), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n600), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n339), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n734), .A2(new_n741), .A3(new_n471), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n734), .B2(new_n723), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n742), .B2(new_n743), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n734), .A2(new_n672), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT114), .B(G78gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  INV_X1    g549(.A(new_n621), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n702), .A2(new_n751), .A3(new_n681), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n698), .A2(new_n657), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G85gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n702), .A2(new_n751), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n584), .B(new_n755), .C1(new_n690), .C2(new_n491), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n483), .A2(new_n492), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n759), .A3(new_n584), .A4(new_n755), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n489), .A2(G85gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n757), .A2(new_n760), .A3(new_n654), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n762), .ZN(G1336gat));
  NAND4_X1  g562(.A1(new_n696), .A2(new_n339), .A3(new_n697), .A4(new_n752), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n367), .A2(G92gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n757), .A2(new_n760), .A3(new_n654), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n770), .A3(KEYINPUT52), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n765), .B(new_n769), .C1(new_n766), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n698), .A2(new_n723), .A3(new_n752), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G99gat), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n669), .A2(G99gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n760), .A3(new_n654), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1338gat));
  NAND4_X1  g578(.A1(new_n696), .A2(new_n672), .A3(new_n697), .A4(new_n752), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G106gat), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n398), .A2(G106gat), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n757), .A2(new_n760), .A3(new_n654), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n642), .B2(new_n645), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n637), .A2(new_n641), .A3(new_n644), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT54), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n626), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n610), .A2(new_n611), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n645), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n647), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n642), .A2(KEYINPUT107), .A3(new_n645), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n789), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(KEYINPUT117), .A3(new_n627), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n795), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n652), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n793), .A2(new_n794), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n805), .A2(KEYINPUT117), .A3(new_n627), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT117), .B1(new_n805), .B2(new_n627), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n702), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n529), .A2(new_n530), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n523), .B1(new_n519), .B2(new_n522), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n539), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n547), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n654), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n584), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n815), .A2(new_n584), .A3(new_n820), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n621), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n655), .A2(new_n703), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n657), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n471), .A2(new_n398), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n828), .A2(new_n339), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n702), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n672), .B1(new_n825), .B2(new_n826), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n669), .A2(new_n489), .A3(new_n339), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n223), .B1(new_n547), .B2(new_n541), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  NOR3_X1   g636(.A1(new_n834), .A2(new_n220), .A3(new_n681), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n830), .A2(new_n654), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n220), .ZN(G1341gat));
  NOR3_X1   g639(.A1(new_n834), .A2(new_n230), .A3(new_n621), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT118), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n830), .A2(new_n751), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(G127gat), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n848), .A3(new_n584), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n834), .B2(new_n683), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n828), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n827), .A2(KEYINPUT123), .A3(new_n657), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n667), .A2(new_n672), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n339), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n680), .A2(new_n208), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n666), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n489), .A2(new_n339), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n398), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n812), .A2(KEYINPUT120), .A3(new_n813), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n809), .B(KEYINPUT55), .C1(new_n810), .C2(new_n811), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n680), .A2(new_n653), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n821), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n870), .A2(new_n808), .A3(new_n680), .A4(new_n871), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n821), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n584), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n823), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n821), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT121), .B1(new_n878), .B2(new_n821), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n683), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT122), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n621), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n868), .B1(new_n887), .B2(new_n826), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n827), .B2(new_n672), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n702), .B(new_n865), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n861), .B1(new_n890), .B2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n824), .B1(new_n885), .B2(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n880), .A2(new_n881), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n751), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n826), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n867), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n889), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n864), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n208), .B1(new_n899), .B2(new_n680), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n892), .B1(new_n901), .B2(new_n859), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n891), .A2(new_n892), .B1(new_n900), .B2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(new_n901), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n210), .A3(new_n654), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n899), .B2(new_n654), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n827), .A2(new_n672), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n751), .B1(new_n885), .B2(new_n823), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n623), .A2(new_n680), .A3(new_n654), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n866), .B(new_n672), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n654), .A3(new_n865), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n905), .B1(new_n908), .B2(new_n915), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n904), .A2(new_n204), .A3(new_n751), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n899), .A2(new_n751), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n204), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n904), .B2(new_n584), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n683), .A2(new_n205), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n899), .B2(new_n921), .ZN(G1347gat));
  AOI21_X1  g721(.A(new_n657), .B1(new_n825), .B2(new_n826), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n829), .A2(new_n367), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n702), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n489), .A2(new_n339), .A3(new_n471), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n832), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n300), .B1(new_n547), .B2(new_n541), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n925), .A2(new_n654), .ZN(new_n933));
  INV_X1    g732(.A(G176gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n929), .A2(new_n299), .A3(new_n681), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(G1349gat));
  NOR2_X1   g737(.A1(new_n621), .A2(new_n287), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G183gat), .B1(new_n929), .B2(new_n621), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n940), .B(new_n941), .C1(KEYINPUT126), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT127), .Z(new_n945));
  XNOR2_X1  g744(.A(new_n943), .B(new_n945), .ZN(G1350gat));
  INV_X1    g745(.A(G190gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n947), .A3(new_n584), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n929), .B2(new_n683), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  AND4_X1   g751(.A1(new_n339), .A2(new_n923), .A3(new_n672), .A4(new_n667), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n702), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n910), .A2(new_n913), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n723), .A2(new_n657), .A3(new_n367), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n680), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  OAI21_X1  g759(.A(G204gat), .B1(new_n957), .B2(new_n681), .ZN(new_n961));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n953), .A2(new_n962), .A3(new_n654), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n953), .A2(new_n276), .A3(new_n751), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n910), .A2(new_n751), .A3(new_n913), .A4(new_n956), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n953), .B2(new_n584), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n683), .A2(new_n275), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n958), .B2(new_n973), .ZN(G1355gat));
endmodule


