//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT81), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT31), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208));
  AND2_X1   g007(.A1(G228gat), .A2(G233gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n215), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT77), .B1(new_n215), .B2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n214), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n210), .B(new_n213), .C1(new_n222), .C2(KEYINPUT2), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  INV_X1    g026(.A(G211gat), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n231), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n225), .B1(new_n236), .B2(KEYINPUT82), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n231), .B(new_n232), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n224), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n243), .B2(KEYINPUT29), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n209), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n247));
  INV_X1    g046(.A(new_n224), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n247), .B(new_n209), .C1(new_n236), .C2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n208), .B(G22gat), .C1(new_n245), .C2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n245), .A2(new_n250), .ZN(new_n252));
  INV_X1    g051(.A(G22gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT84), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(G22gat), .B1(new_n245), .B2(new_n250), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n207), .B(new_n251), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258));
  INV_X1    g057(.A(new_n250), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(new_n239), .B2(new_n240), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n240), .B2(new_n239), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n246), .B1(new_n261), .B2(new_n224), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n253), .B(new_n259), .C1(new_n262), .C2(new_n209), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n255), .ZN(new_n264));
  INV_X1    g063(.A(new_n207), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI211_X1 g065(.A(KEYINPUT83), .B(new_n207), .C1(new_n263), .C2(new_n255), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n257), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT27), .B(G183gat), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT28), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  OR3_X1    g072(.A1(new_n273), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT27), .B1(new_n273), .B2(KEYINPUT69), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n270), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(KEYINPUT26), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n280), .A2(new_n281), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n286), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  OR2_X1    g093(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n295));
  INV_X1    g094(.A(new_n289), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n296), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n291), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n293), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT25), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT66), .B(G176gat), .Z(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(new_n291), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT25), .B1(new_n304), .B2(new_n282), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n294), .B1(new_n296), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n289), .A2(KEYINPUT64), .A3(new_n306), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n300), .A2(new_n286), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n308), .A2(new_n314), .A3(new_n309), .A4(new_n310), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n305), .A2(new_n312), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n290), .A2(new_n302), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT71), .A3(G134gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT72), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n320), .A2(new_n328), .A3(new_n322), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G227gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n290), .A2(new_n302), .A3(new_n316), .ZN(new_n337));
  INV_X1    g136(.A(new_n331), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n327), .B2(new_n329), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n343));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G71gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G99gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n341), .A2(new_n349), .A3(KEYINPUT32), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(new_n336), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n336), .B(new_n352), .C1(new_n333), .C2(new_n340), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n341), .B(KEYINPUT32), .C1(new_n347), .C2(new_n346), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n351), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n351), .A2(new_n359), .ZN(new_n361));
  INV_X1    g160(.A(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n268), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n202), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n332), .A2(new_n224), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n248), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n339), .A2(new_n243), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(new_n247), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n374), .B2(new_n247), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n339), .A2(new_n379), .A3(new_n248), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n379), .A4(new_n248), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n373), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G57gat), .ZN(new_n389));
  INV_X1    g188(.A(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n247), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT78), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n247), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n383), .A2(new_n380), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n367), .A3(new_n371), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT80), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n386), .B2(new_n397), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n403), .A3(new_n397), .A4(new_n391), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n399), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(KEYINPUT6), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n337), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n317), .A2(KEYINPUT29), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n234), .B(new_n409), .C1(new_n410), .C2(new_n408), .ZN(new_n411));
  INV_X1    g210(.A(new_n409), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n337), .B2(new_n235), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n238), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT75), .ZN(new_n416));
  INV_X1    g215(.A(G64gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G92gat), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT30), .A4(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(new_n414), .ZN(new_n422));
  INV_X1    g221(.A(new_n419), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n411), .A2(new_n414), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n364), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n366), .A2(new_n407), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n360), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n358), .B1(new_n351), .B2(new_n359), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT88), .A3(new_n268), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n268), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n407), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n202), .B(new_n435), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n405), .B2(new_n406), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n442), .A2(new_n268), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n370), .B2(new_n372), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT86), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(KEYINPUT39), .C1(new_n370), .C2(new_n372), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n393), .A2(new_n394), .B1(new_n383), .B2(new_n380), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n447), .C1(new_n448), .C2(new_n371), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n395), .A2(new_n396), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT85), .B(KEYINPUT39), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n372), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT40), .A4(new_n391), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n452), .A3(new_n391), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n429), .A2(new_n401), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n422), .A2(new_n423), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n422), .A2(KEYINPUT37), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n411), .A2(new_n414), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n423), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT38), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n423), .A3(new_n461), .A4(new_n459), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n457), .B(new_n268), .C1(new_n407), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n432), .B2(new_n433), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n443), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n441), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G120gat), .B(G148gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(new_n283), .ZN(new_n479));
  INV_X1    g278(.A(G204gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G57gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G64gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n417), .A2(G57gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT96), .ZN(new_n491));
  INV_X1    g290(.A(new_n485), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G71gat), .B(G78gat), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n486), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n486), .B2(new_n493), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT102), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G99gat), .ZN(new_n502));
  INV_X1    g301(.A(G106gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT102), .ZN(new_n505));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT7), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(G85gat), .A3(G92gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G92gat), .ZN(new_n514));
  AOI22_X1  g313(.A1(KEYINPUT8), .A2(new_n506), .B1(new_n390), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n507), .A3(new_n513), .A4(new_n515), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT104), .B1(new_n498), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT104), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(new_n522), .C1(new_n496), .C2(new_n497), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n484), .A2(KEYINPUT96), .A3(new_n485), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT95), .B1(new_n490), .B2(new_n492), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n494), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n486), .A2(new_n493), .A3(new_n495), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n518), .A3(new_n517), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT105), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT105), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n519), .A2(new_n532), .A3(new_n528), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n524), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n530), .A2(KEYINPUT106), .A3(new_n525), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT106), .B1(new_n530), .B2(new_n525), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT109), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n534), .ZN(new_n543));
  INV_X1    g342(.A(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n482), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT108), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT107), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n520), .A2(new_n523), .B1(new_n531), .B2(new_n533), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n550), .A2(new_n525), .B1(new_n537), .B2(new_n536), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n551), .B2(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n539), .A2(KEYINPUT107), .A3(new_n540), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n545), .A2(new_n482), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n548), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT108), .B(new_n555), .C1(new_n552), .C2(new_n553), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n547), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT110), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT107), .B1(new_n539), .B2(new_n540), .ZN(new_n561));
  AOI211_X1 g360(.A(new_n549), .B(new_n544), .C1(new_n535), .C2(new_n538), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT108), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n548), .A3(new_n556), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT110), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n547), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(G1gat), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT90), .B(G29gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G36gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(G29gat), .B2(G36gat), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n580), .A2(G29gat), .A3(G36gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT91), .B(G50gat), .ZN(new_n584));
  INV_X1    g383(.A(G43gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT15), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n204), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT92), .ZN(new_n591));
  NOR2_X1   g390(.A1(G43gat), .A2(G50gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT15), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n583), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n583), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n586), .A2(new_n597), .A3(new_n587), .A4(new_n589), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n577), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n596), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n593), .B1(new_n603), .B2(new_n583), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT93), .A4(KEYINPUT17), .ZN(new_n605));
  OR2_X1    g404(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n606), .B(new_n607), .C1(new_n594), .C2(new_n599), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n600), .B1(new_n609), .B2(new_n577), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n611), .B(KEYINPUT13), .Z(new_n615));
  NOR2_X1   g414(.A1(new_n594), .A2(new_n599), .ZN(new_n616));
  INV_X1    g415(.A(new_n577), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n615), .B1(new_n618), .B2(new_n600), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT94), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n621), .B(new_n615), .C1(new_n618), .C2(new_n600), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n614), .A2(new_n623), .A3(new_n633), .A4(new_n624), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n569), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n609), .A2(new_n521), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n519), .ZN(new_n639));
  NAND3_X1  g438(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G190gat), .B(G218gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(G134gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G162gat), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n643), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(KEYINPUT103), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n644), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n617), .B1(KEYINPUT21), .B2(new_n498), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n498), .A2(KEYINPUT21), .ZN(new_n655));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT97), .ZN(new_n660));
  XOR2_X1   g459(.A(G183gat), .B(G211gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n658), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n477), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n438), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n573), .A2(new_n572), .ZN(new_n673));
  NAND2_X1  g472(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n674));
  AND4_X1   g473(.A1(new_n429), .A2(new_n670), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n572), .B1(new_n670), .B2(new_n429), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n675), .ZN(G1325gat));
  AOI21_X1  g477(.A(G15gat), .B1(new_n670), .B2(new_n434), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n472), .A2(new_n474), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n670), .B2(new_n681), .ZN(G1326gat));
  INV_X1    g481(.A(new_n268), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n670), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n687), .A3(new_n683), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n685), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n253), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(G22gat), .A3(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n477), .A2(new_n651), .ZN(new_n696));
  INV_X1    g495(.A(new_n667), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n637), .A2(new_n697), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n696), .A2(new_n407), .A3(new_n578), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  AND4_X1   g500(.A1(new_n405), .A2(new_n466), .A3(new_n469), .A4(new_n406), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n456), .A2(new_n401), .A3(new_n453), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n268), .B1(new_n703), .B2(new_n436), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n702), .A2(new_n704), .B1(new_n442), .B2(new_n268), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT112), .B1(new_n705), .B2(new_n680), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n443), .A2(new_n471), .A3(new_n707), .A4(new_n475), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n440), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n701), .B1(new_n709), .B2(new_n652), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n477), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n637), .A4(new_n697), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n578), .B1(new_n712), .B2(new_n407), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n700), .A2(new_n713), .ZN(G1328gat));
  NOR4_X1   g513(.A1(new_n696), .A2(G36gat), .A3(new_n436), .A4(new_n698), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n436), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  OAI21_X1  g517(.A(G43gat), .B1(new_n712), .B2(new_n475), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n696), .A2(new_n698), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n585), .A3(new_n434), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n584), .A3(new_n683), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n712), .A2(new_n268), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n584), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n726), .B(new_n728), .ZN(G1331gat));
  INV_X1    g528(.A(new_n569), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n668), .A2(new_n635), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n709), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n438), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  INV_X1    g534(.A(new_n733), .ZN(new_n736));
  AOI211_X1 g535(.A(new_n436), .B(new_n736), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n733), .A2(G71gat), .A3(new_n680), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n733), .A2(new_n434), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G71gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n683), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n667), .A2(new_n635), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n710), .A2(new_n711), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT114), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n710), .A2(new_n711), .A3(new_n751), .A4(new_n748), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n407), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n706), .A2(new_n708), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n652), .B1(new_n754), .B2(new_n441), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT51), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NOR4_X1   g556(.A1(new_n709), .A2(new_n757), .A3(new_n652), .A4(new_n747), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n569), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n438), .A2(new_n390), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n753), .A2(new_n390), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n752), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n514), .B1(new_n762), .B2(new_n429), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n514), .B(new_n569), .C1(new_n756), .C2(new_n758), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n436), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n749), .B2(new_n436), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1337gat));
  AOI21_X1  g569(.A(new_n475), .B1(new_n750), .B2(new_n752), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n434), .A2(new_n502), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n771), .A2(new_n502), .B1(new_n759), .B2(new_n772), .ZN(G1338gat));
  AOI21_X1  g572(.A(new_n503), .B1(new_n762), .B2(new_n683), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n569), .A2(new_n683), .A3(new_n503), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT115), .Z(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n756), .B2(new_n758), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT116), .B(new_n776), .C1(new_n756), .C2(new_n758), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n749), .B2(new_n268), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n756), .A2(new_n758), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n775), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n407), .A2(new_n429), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n610), .A2(new_n611), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n618), .A2(new_n600), .A3(new_n615), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n630), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n634), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT117), .ZN(new_n793));
  OAI221_X1 g592(.A(KEYINPUT54), .B1(new_n539), .B2(new_n541), .C1(new_n561), .C2(new_n562), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n481), .B1(new_n542), .B2(KEYINPUT54), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n566), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n539), .A2(new_n541), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n552), .B2(new_n553), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n795), .B1(new_n800), .B2(KEYINPUT54), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n801), .A2(KEYINPUT55), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n793), .A2(new_n651), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n567), .B1(new_n566), .B2(new_n547), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT110), .B(new_n546), .C1(new_n564), .C2(new_n565), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n792), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n798), .A2(new_n635), .A3(new_n802), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n651), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n697), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n731), .A2(new_n730), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n683), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n434), .B(new_n788), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n635), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G113gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n810), .A2(new_n811), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n438), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n437), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n823), .A2(G113gat), .A3(new_n636), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n824), .ZN(G1340gat));
  NAND3_X1  g624(.A1(new_n816), .A2(new_n817), .A3(new_n569), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G120gat), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n823), .A2(G120gat), .A3(new_n730), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1341gat));
  NAND4_X1  g628(.A1(new_n816), .A2(new_n817), .A3(G127gat), .A4(new_n667), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n321), .B1(new_n823), .B2(new_n697), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n651), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G134gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n823), .A2(G134gat), .A3(new_n652), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1343gat));
  AND2_X1   g636(.A1(new_n475), .A2(new_n788), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n683), .A2(KEYINPUT57), .ZN(new_n839));
  INV_X1    g638(.A(new_n792), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n560), .B2(new_n568), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n635), .B1(KEYINPUT55), .B2(new_n801), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n797), .A2(new_n566), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT120), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n807), .A2(new_n846), .A3(new_n808), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n652), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT121), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(new_n847), .A3(new_n850), .A4(new_n652), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n803), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n697), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n839), .B1(new_n853), .B2(new_n811), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n820), .B2(new_n683), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n635), .B(new_n838), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n821), .A2(KEYINPUT122), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n268), .A3(new_n680), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n429), .B1(new_n821), .B2(KEYINPUT122), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n219), .A3(new_n635), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n861), .A3(new_n863), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1344gat));
  AND2_X1   g666(.A1(new_n859), .A2(new_n860), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n215), .A3(new_n569), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n838), .B1(new_n854), .B2(new_n855), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n730), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n215), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n667), .B1(new_n848), .B2(new_n803), .ZN(new_n874));
  INV_X1    g673(.A(new_n811), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n820), .A2(new_n683), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n877), .A2(new_n683), .B1(KEYINPUT57), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n569), .A3(new_n838), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n870), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n869), .B1(new_n873), .B2(new_n881), .ZN(G1345gat));
  AOI21_X1  g681(.A(G155gat), .B1(new_n868), .B2(new_n667), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n871), .A2(new_n211), .A3(new_n697), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n212), .A3(new_n651), .ZN(new_n886));
  OAI21_X1  g685(.A(G162gat), .B1(new_n871), .B2(new_n652), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n438), .A2(new_n436), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n434), .B(new_n889), .C1(new_n813), .C2(new_n814), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n636), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n438), .B1(new_n810), .B2(new_n811), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n268), .A2(new_n892), .A3(new_n434), .A4(new_n429), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n282), .A3(new_n635), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n893), .B2(new_n569), .ZN(new_n896));
  INV_X1    g695(.A(new_n890), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n569), .A2(new_n303), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n890), .B2(new_n697), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n269), .A3(new_n667), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g702(.A1(new_n890), .A2(new_n652), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n270), .ZN(new_n905));
  NAND2_X1  g704(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n270), .A3(new_n651), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n907), .B(new_n908), .C1(new_n904), .C2(new_n270), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G1351gat));
  NAND3_X1  g712(.A1(new_n475), .A2(new_n683), .A3(new_n429), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n635), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n889), .A2(new_n475), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n879), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n635), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(new_n920), .ZN(G1352gat));
  NOR3_X1   g724(.A1(new_n918), .A2(G204gat), .A3(new_n730), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(KEYINPUT126), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n879), .A2(new_n569), .A3(new_n922), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n930), .B(new_n931), .C1(new_n480), .C2(new_n932), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n228), .A3(new_n667), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n879), .A2(new_n667), .A3(new_n922), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n919), .B2(new_n651), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n651), .A2(G218gat), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT127), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n923), .B2(new_n941), .ZN(G1355gat));
endmodule


