//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1207,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n212), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT64), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n215), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g0043(.A1(G68), .A2(G77), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT76), .ZN(new_n250));
  INV_X1    g0050(.A(G58), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n201), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G58), .A2(G68), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G159), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT16), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT74), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(G20), .B1(new_n262), .B2(new_n264), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT74), .B1(new_n271), .B2(KEYINPUT7), .ZN(new_n272));
  OAI21_X1  g0072(.A(G68), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT75), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT75), .B(G68), .C1(new_n270), .C2(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n260), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n263), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT7), .B(new_n210), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G68), .ZN(new_n282));
  INV_X1    g0082(.A(new_n257), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT16), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n285), .A2(new_n226), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n277), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n289), .A2(new_n251), .A3(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n286), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n209), .B2(G20), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n294), .B1(new_n296), .B2(new_n292), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n250), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n276), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT74), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n269), .A3(new_n266), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT75), .B1(new_n303), .B2(G68), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n259), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n284), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n295), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT76), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n268), .A2(G226), .A3(G1698), .ZN(new_n309));
  INV_X1    g0109(.A(G1698), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G41), .ZN(new_n316));
  INV_X1    g0116(.A(G45), .ZN(new_n317));
  AOI21_X1  g0117(.A(G1), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT68), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G41), .A2(G45), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(G1), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G274), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n314), .A2(new_n318), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n323), .A2(new_n325), .B1(new_n326), .B2(G232), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n315), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(G169), .B1(new_n315), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT77), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n315), .A2(new_n327), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n315), .A2(new_n327), .A3(new_n328), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n299), .A2(new_n308), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT18), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n299), .A2(new_n341), .A3(new_n308), .A4(new_n338), .ZN(new_n342));
  INV_X1    g0142(.A(G200), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(G190), .B2(new_n332), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n307), .A2(new_n345), .A3(new_n297), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT17), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n340), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n323), .A2(new_n325), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G226), .B2(new_n326), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n268), .A2(G222), .A3(new_n310), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n268), .A2(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G223), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n351), .B1(new_n202), .B2(new_n268), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n314), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(G200), .B2(new_n356), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n210), .A2(G33), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n292), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G50), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n251), .A3(new_n201), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n286), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n296), .A2(G50), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G50), .B2(new_n293), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(KEYINPUT9), .B1(KEYINPUT70), .B2(KEYINPUT10), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(KEYINPUT9), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n359), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n368), .B1(new_n333), .B2(new_n356), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G179), .B2(new_n356), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n296), .A2(G68), .ZN(new_n378));
  XOR2_X1   g0178(.A(new_n378), .B(KEYINPUT71), .Z(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT72), .B1(new_n293), .B2(G68), .ZN(new_n380));
  XOR2_X1   g0180(.A(new_n380), .B(KEYINPUT12), .Z(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n255), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n362), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n360), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n295), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g0186(.A(new_n386), .B(KEYINPUT11), .Z(new_n387));
  NOR2_X1   g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n268), .A2(G226), .A3(new_n310), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n314), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n323), .A2(new_n325), .B1(new_n326), .B2(G238), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G179), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n407), .A3(G169), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n389), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(G200), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n397), .A2(G190), .A3(new_n399), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n388), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n296), .A2(G77), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G77), .B2(new_n293), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G20), .A2(G77), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n417), .B1(new_n288), .B2(new_n383), .C1(new_n360), .C2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n295), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n349), .B1(G244), .B2(new_n326), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n268), .A2(G232), .A3(new_n310), .ZN(new_n422));
  INV_X1    g0222(.A(G238), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n206), .B2(new_n268), .C1(new_n352), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n314), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n420), .B1(new_n426), .B2(new_n333), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n328), .A3(new_n425), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n420), .C1(new_n357), .C2(new_n426), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n348), .A2(new_n377), .A3(new_n414), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT6), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n434), .A2(new_n205), .A3(G107), .ZN(new_n435));
  XNOR2_X1  g0235(.A(G97), .B(G107), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n437), .A2(new_n210), .B1(new_n202), .B2(new_n383), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n206), .B1(new_n269), .B2(new_n280), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n295), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n293), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n209), .A2(G33), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n286), .A2(new_n293), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n443), .B2(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT78), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n268), .A2(G244), .A3(new_n310), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n449), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n268), .A2(new_n451), .A3(G244), .A4(new_n310), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n314), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  OAI211_X1 g0257(.A(G1), .B(G13), .C1(new_n261), .C2(new_n316), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n209), .A2(G45), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AND4_X1   g0260(.A1(G274), .A2(new_n457), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n314), .B1(new_n460), .B2(new_n457), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(G257), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G200), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT78), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n440), .A2(new_n466), .A3(new_n444), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n456), .A2(G190), .A3(new_n463), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n446), .A2(new_n465), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n456), .A2(G179), .A3(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n333), .B1(new_n456), .B2(new_n463), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n445), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT80), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n458), .A2(G274), .A3(new_n460), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n458), .A2(G250), .A3(new_n459), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n268), .A2(G244), .A3(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n262), .A2(new_n264), .A3(G238), .A4(new_n310), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n328), .B(new_n478), .C1(new_n314), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n314), .ZN(new_n484));
  INV_X1    g0284(.A(new_n478), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n333), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n475), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(G179), .A3(new_n485), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n478), .B1(new_n482), .B2(new_n314), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(KEYINPUT80), .C1(new_n333), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n268), .A2(new_n210), .A3(G68), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n210), .B1(new_n392), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(G87), .B2(new_n207), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n360), .B2(new_n205), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n293), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n496), .A2(new_n295), .B1(new_n497), .B2(new_n418), .ZN(new_n498));
  INV_X1    g0298(.A(new_n418), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n443), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n487), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n484), .A2(new_n485), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n357), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n489), .A2(new_n343), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n443), .A2(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  OR3_X1    g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n474), .A2(new_n510), .A3(KEYINPUT81), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n469), .A2(new_n473), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n206), .A3(G20), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n268), .A2(new_n210), .A3(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n268), .A2(new_n525), .A3(new_n210), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n522), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n295), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT25), .B1(new_n497), .B2(new_n206), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n497), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n443), .B2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n262), .A2(new_n264), .A3(G250), .A4(new_n310), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n314), .B1(G264), .B2(new_n462), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n325), .A2(new_n460), .A3(new_n457), .ZN(new_n542));
  AOI21_X1  g0342(.A(G169), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n541), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n461), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n543), .B1(new_n545), .B2(new_n328), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n541), .A2(new_n357), .A3(new_n542), .ZN(new_n550));
  AOI21_X1  g0350(.A(G200), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT85), .B(G200), .C1(new_n541), .C2(new_n542), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n531), .B(new_n535), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n536), .A2(new_n546), .A3(KEYINPUT84), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n443), .A2(G116), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n497), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n285), .A2(new_n226), .B1(G20), .B2(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n453), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT20), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n558), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n461), .B1(G270), .B2(new_n462), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n268), .A2(G257), .A3(new_n310), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n268), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n314), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n567), .A2(new_n572), .A3(G179), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(G169), .A3(new_n565), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT82), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n565), .B1(new_n573), .B2(G200), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n357), .B2(new_n573), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n557), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n433), .A2(new_n515), .A3(new_n585), .ZN(G372));
  NAND2_X1  g0386(.A1(new_n410), .A2(new_n429), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n347), .A3(new_n413), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n331), .A2(new_n337), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n307), .B2(new_n297), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n374), .A3(new_n373), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(new_n376), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT86), .B1(new_n483), .B2(new_n486), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT86), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n488), .B(new_n597), .C1(new_n333), .C2(new_n489), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n595), .B1(new_n599), .B2(new_n501), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n600), .A2(new_n473), .A3(new_n469), .A4(new_n555), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n580), .A2(new_n581), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n603), .B2(new_n547), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT26), .B1(new_n509), .B2(new_n473), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n501), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n464), .A2(G169), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n446), .A2(new_n467), .B1(new_n607), .B2(new_n470), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT26), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n606), .A2(new_n608), .A3(new_n609), .A4(new_n508), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n605), .A2(new_n610), .A3(new_n606), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n433), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n594), .A2(new_n612), .ZN(G369));
  NAND3_X1  g0413(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(KEYINPUT27), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(KEYINPUT27), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(G213), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(G343), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(G343), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n602), .A2(new_n565), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n566), .A2(new_n623), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n584), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(G330), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n623), .B1(new_n531), .B2(new_n535), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n557), .A2(new_n629), .B1(new_n547), .B2(new_n623), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n536), .A2(new_n546), .A3(new_n623), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n603), .A2(new_n624), .ZN(new_n633));
  INV_X1    g0433(.A(new_n557), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(G399));
  INV_X1    g0436(.A(new_n213), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(G41), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G1), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n225), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(new_n639), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT28), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n605), .A2(new_n610), .A3(new_n606), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n555), .A2(new_n473), .A3(new_n469), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n580), .A2(new_n581), .A3(new_n547), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n600), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n624), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT88), .B1(new_n649), .B2(KEYINPUT29), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n623), .B1(new_n604), .B2(new_n611), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT29), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n536), .A2(new_n546), .A3(KEYINPUT84), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT84), .B1(new_n536), .B2(new_n546), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n601), .B1(new_n603), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n607), .A2(new_n470), .B1(new_n440), .B2(new_n444), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(new_n502), .A3(new_n609), .A4(new_n508), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n446), .A2(new_n467), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n607), .A2(new_n470), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n596), .A2(new_n598), .B1(new_n498), .B2(new_n500), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n665), .A3(new_n595), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n606), .B(new_n661), .C1(new_n666), .C2(new_n609), .ZN(new_n667));
  OAI211_X1 g0467(.A(KEYINPUT29), .B(new_n623), .C1(new_n659), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT89), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n661), .A2(new_n606), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n600), .A2(new_n608), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(KEYINPUT26), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n549), .A2(new_n556), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n646), .B(new_n600), .C1(new_n673), .C2(new_n602), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT29), .A4(new_n623), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n655), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n515), .A2(new_n585), .A3(new_n623), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n456), .A2(new_n463), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n544), .A2(new_n503), .ZN(new_n682));
  INV_X1    g0482(.A(new_n575), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n573), .A2(new_n328), .A3(new_n503), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n687), .B(new_n464), .C1(new_n461), .C2(new_n544), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(KEYINPUT30), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n624), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n680), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n679), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n644), .B1(new_n697), .B2(G1), .ZN(G364));
  INV_X1    g0498(.A(G13), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G20), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n209), .B1(new_n700), .B2(G45), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n638), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n628), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G330), .B2(new_n627), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n213), .A2(new_n268), .ZN(new_n706));
  INV_X1    g0506(.A(G355), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(G116), .B2(new_n213), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n248), .A2(G45), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n268), .B(new_n637), .C1(new_n317), .C2(new_n225), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n226), .B1(G20), .B2(new_n333), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n703), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n210), .A2(new_n357), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n343), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n328), .A2(G200), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n210), .A2(G190), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(new_n726), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n728), .A2(new_n251), .B1(new_n731), .B2(new_n202), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT90), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n725), .A2(G87), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n720), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n268), .B1(new_n735), .B2(new_n206), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G179), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n740), .B2(KEYINPUT32), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n734), .B(new_n741), .C1(new_n733), .C2(new_n732), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n210), .A2(new_n328), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n210), .B1(new_n737), .B2(G190), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n362), .B1(new_n745), .B2(new_n205), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(new_n357), .A3(G200), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n740), .A2(KEYINPUT32), .B1(new_n201), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n742), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  OAI22_X1  g0554(.A1(new_n728), .A2(new_n753), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  AOI22_X1  g0556(.A1(G329), .A2(new_n739), .B1(new_n730), .B2(G311), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n265), .C1(new_n758), .C2(new_n735), .ZN(new_n759));
  INV_X1    g0559(.A(G326), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n744), .A2(new_n760), .B1(new_n745), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n756), .B(new_n763), .C1(new_n570), .C2(new_n724), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n751), .A2(new_n752), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n718), .B1(new_n765), .B2(new_n715), .ZN(new_n766));
  INV_X1    g0566(.A(new_n714), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n627), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n705), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(G396));
  OAI21_X1  g0570(.A(new_n431), .B1(new_n420), .B2(new_n623), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n429), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n427), .A2(new_n428), .A3(new_n623), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n649), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n696), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(KEYINPUT96), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(KEYINPUT96), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n777), .A2(new_n778), .A3(new_n703), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n696), .A2(new_n775), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n779), .B2(KEYINPUT97), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n703), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n715), .A2(new_n712), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G77), .ZN(new_n788));
  INV_X1    g0588(.A(new_n747), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G283), .B1(new_n730), .B2(G116), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  INV_X1    g0591(.A(new_n744), .ZN(new_n792));
  INV_X1    g0592(.A(new_n745), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G303), .B1(new_n793), .B2(G97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n735), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G87), .A2(new_n795), .B1(new_n739), .B2(G311), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n268), .B1(new_n727), .B2(G294), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n791), .B(new_n798), .C1(new_n206), .C2(new_n724), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G143), .A2(new_n727), .B1(new_n730), .B2(G159), .ZN(new_n800));
  INV_X1    g0600(.A(G150), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n747), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G137), .B2(new_n792), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT34), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n268), .B1(new_n735), .B2(new_n201), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G132), .B2(new_n739), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n251), .B2(new_n745), .C1(new_n362), .C2(new_n724), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n799), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT95), .ZN(new_n809));
  INV_X1    g0609(.A(new_n715), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n808), .B2(KEYINPUT95), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n785), .B(new_n788), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n774), .A2(new_n712), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n784), .A2(new_n814), .ZN(G384));
  OAI21_X1  g0615(.A(new_n283), .B1(new_n300), .B2(new_n304), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n258), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n275), .A2(new_n276), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n286), .B1(new_n818), .B2(new_n259), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n298), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n346), .B1(new_n820), .B2(new_n617), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n589), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT37), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n299), .A2(new_n308), .A3(new_n618), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n307), .A2(new_n297), .A3(new_n345), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n339), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n820), .A2(new_n617), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n348), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n831), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT38), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT102), .B1(new_n828), .B2(new_n590), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n338), .B1(new_n287), .B2(new_n298), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT102), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n346), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n827), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n339), .A2(new_n829), .ZN(new_n844));
  AOI22_X1  g0644(.A1(KEYINPUT37), .A2(new_n843), .B1(new_n844), .B2(new_n827), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n827), .B1(new_n591), .B2(new_n347), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n831), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT39), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n410), .A2(new_n624), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n837), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n834), .A2(new_n835), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n773), .B1(new_n651), .B2(new_n774), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n388), .A2(new_n623), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n414), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n410), .B(new_n413), .C1(new_n388), .C2(new_n623), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n853), .A2(new_n859), .B1(new_n591), .B2(new_n618), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n655), .A2(new_n678), .A3(new_n433), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n594), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n861), .B(new_n863), .Z(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n691), .B2(new_n692), .ZN(new_n867));
  AOI211_X1 g0667(.A(KEYINPUT104), .B(KEYINPUT31), .C1(new_n690), .C2(new_n624), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n680), .A3(new_n694), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n774), .B1(new_n856), .B2(new_n857), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n865), .B1(new_n853), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n830), .ZN(new_n876));
  INV_X1    g0676(.A(new_n846), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n874), .B(KEYINPUT40), .C1(new_n834), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n433), .A2(new_n870), .ZN(new_n881));
  OAI21_X1  g0681(.A(G330), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n864), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n864), .A2(new_n883), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(new_n885), .C1(new_n209), .C2(new_n700), .ZN(new_n886));
  INV_X1    g0686(.A(new_n437), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n887), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n227), .A4(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n642), .A2(new_n202), .A3(new_n252), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n201), .A2(G50), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT100), .Z(new_n897));
  NOR3_X1   g0697(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n699), .A2(G1), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n886), .B(new_n891), .C1(new_n898), .C2(new_n899), .ZN(G367));
  INV_X1    g0700(.A(new_n697), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n635), .A2(new_n632), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n623), .B1(new_n446), .B2(new_n467), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n513), .A2(new_n903), .B1(new_n664), .B2(new_n623), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT44), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(KEYINPUT106), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n635), .A2(new_n632), .A3(new_n904), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT45), .Z(new_n911));
  AND3_X1   g0711(.A1(new_n909), .A2(new_n911), .A3(new_n631), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n631), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n635), .B1(new_n630), .B2(new_n633), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(new_n628), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n697), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n909), .A2(new_n911), .ZN(new_n919));
  INV_X1    g0719(.A(new_n631), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n909), .A2(new_n911), .A3(new_n631), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n697), .A2(new_n917), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT107), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n901), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n638), .B(KEYINPUT41), .Z(new_n927));
  OAI21_X1  g0727(.A(new_n701), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n633), .A2(new_n634), .A3(new_n904), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT42), .Z(new_n930));
  AND2_X1   g0730(.A1(new_n904), .A2(new_n673), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n623), .B1(new_n931), .B2(new_n660), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n507), .A2(new_n624), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n600), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n665), .A2(new_n507), .A3(new_n624), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT43), .B1(new_n937), .B2(KEYINPUT105), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(KEYINPUT105), .B2(new_n937), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n933), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n920), .A2(new_n904), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n942), .B(new_n943), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n928), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n745), .A2(new_n201), .ZN(new_n946));
  INV_X1    g0746(.A(G159), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n268), .B1(new_n947), .B2(new_n747), .C1(new_n728), .C2(new_n801), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(G143), .C2(new_n792), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n795), .A2(G77), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n362), .B2(new_n731), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G137), .B2(new_n739), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n949), .B(new_n952), .C1(new_n251), .C2(new_n724), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT108), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n795), .A2(G97), .B1(new_n727), .B2(G303), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n758), .B2(new_n731), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n268), .B1(new_n739), .B2(G317), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n761), .B2(new_n747), .ZN(new_n958));
  INV_X1    g0758(.A(G311), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n744), .A2(new_n959), .B1(new_n745), .B2(new_n206), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n724), .A2(new_n559), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT46), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n954), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n715), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n716), .B1(new_n213), .B2(new_n418), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n637), .A2(new_n268), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n237), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n785), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n966), .B(new_n970), .C1(new_n767), .C2(new_n937), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n945), .A2(new_n971), .ZN(G387));
  NAND2_X1  g0772(.A1(new_n917), .A2(new_n702), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G317), .A2(new_n727), .B1(new_n730), .B2(G303), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n959), .B2(new_n747), .C1(new_n753), .C2(new_n744), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT48), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n724), .A2(new_n761), .B1(new_n758), .B2(new_n745), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT111), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT112), .Z(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT49), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT49), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n265), .B1(new_n738), .B2(new_n760), .C1(new_n559), .C2(new_n735), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n731), .A2(new_n201), .B1(new_n738), .B2(new_n801), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G50), .B2(new_n727), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n725), .A2(G77), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n745), .A2(new_n418), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n268), .B1(new_n735), .B2(new_n205), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G159), .C2(new_n792), .ZN(new_n990));
  INV_X1    g0790(.A(new_n292), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n789), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n987), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n810), .B1(new_n984), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT113), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n706), .A2(new_n640), .B1(G107), .B2(new_n213), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT109), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n288), .A2(G50), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT50), .Z(new_n999));
  NAND3_X1  g0799(.A1(new_n640), .A2(new_n317), .A3(new_n244), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n968), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n997), .A2(new_n1001), .B1(new_n234), .B2(G45), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n997), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n703), .B1(new_n1004), .B2(new_n717), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT110), .Z(new_n1006));
  OR3_X1    g0806(.A1(new_n994), .A2(new_n995), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n995), .B1(new_n994), .B2(new_n1006), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n630), .C2(new_n767), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n638), .B(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n924), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n697), .A2(new_n917), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n973), .B(new_n1009), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT115), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(G393));
  AND2_X1   g0817(.A1(new_n242), .A2(new_n968), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n716), .B1(new_n205), .B2(new_n213), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n703), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n792), .A2(G317), .B1(new_n727), .B2(G311), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n725), .A2(G283), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n268), .B1(new_n795), .B2(G107), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G322), .A2(new_n739), .B1(new_n730), .B2(G294), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n789), .A2(G303), .B1(new_n793), .B2(G116), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n725), .A2(G68), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n265), .B1(new_n795), .B2(G87), .ZN(new_n1029));
  INV_X1    g0829(.A(G143), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n731), .A2(new_n288), .B1(new_n738), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n745), .A2(new_n202), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G50), .B2(new_n789), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n792), .A2(G150), .B1(new_n727), .B2(G159), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1022), .A2(new_n1027), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1020), .B1(new_n715), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n904), .B2(new_n767), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT116), .B1(new_n912), .B2(new_n913), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT116), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n922), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1041), .B1(new_n1045), .B2(new_n701), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n918), .A2(new_n925), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1010), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(new_n924), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G390));
  OAI21_X1  g0851(.A(new_n712), .B1(new_n837), .B2(new_n849), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n703), .B1(new_n991), .B2(new_n787), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n728), .A2(new_n559), .B1(new_n731), .B2(new_n205), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G294), .B2(new_n739), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n725), .A2(G87), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n268), .B(new_n1033), .C1(G68), .C2(new_n795), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n789), .A2(G107), .B1(new_n792), .B2(G283), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n724), .A2(KEYINPUT53), .A3(new_n801), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT53), .B1(new_n724), .B2(new_n801), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT54), .B(G143), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n789), .A2(G137), .B1(new_n730), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1060), .B(new_n1061), .C1(KEYINPUT121), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(KEYINPUT121), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n265), .B1(new_n795), .B2(G50), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G132), .A2(new_n727), .B1(new_n739), .B2(G125), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n792), .A2(G128), .B1(new_n793), .B2(G159), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1059), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1053), .B1(new_n1072), .B2(new_n715), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1052), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n870), .A2(new_n871), .A3(G330), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n850), .B1(new_n854), .B2(new_n858), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n836), .B1(new_n834), .B2(new_n878), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n831), .A2(new_n833), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n838), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n834), .A2(new_n878), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n773), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n624), .B1(new_n672), .B2(new_n674), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n772), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n858), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n851), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1076), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1077), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n837), .B2(new_n849), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n774), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n695), .A2(G330), .A3(new_n1094), .A4(new_n858), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1074), .B1(new_n1097), .B2(new_n701), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n433), .A2(G330), .A3(new_n870), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n862), .A2(new_n594), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n695), .A2(G330), .A3(new_n1094), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n1087), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n854), .B1(new_n1103), .B2(new_n1076), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n870), .A2(G330), .A3(new_n1094), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1086), .B(new_n1095), .C1(new_n1105), .C2(new_n858), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1101), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1097), .B2(KEYINPUT120), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(KEYINPUT120), .B2(new_n1097), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1090), .A2(new_n1096), .A3(new_n1107), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1090), .A2(new_n1096), .A3(new_n1107), .A4(KEYINPUT118), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1048), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT119), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(KEYINPUT119), .B(new_n1048), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1099), .B1(new_n1116), .B2(new_n1117), .ZN(G378));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1101), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT122), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT57), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n368), .A2(new_n617), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n377), .B(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1128), .A2(new_n873), .A3(G330), .A4(new_n879), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n872), .B1(new_n1080), .B2(new_n848), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n865), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n879), .B(G330), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1127), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n861), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n861), .A3(new_n1129), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1123), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1121), .A2(new_n1122), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1101), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1133), .A2(new_n861), .A3(new_n1129), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n1134), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1123), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT57), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT122), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1138), .A2(new_n1142), .A3(new_n1144), .A4(new_n1010), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n265), .A2(new_n316), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G107), .B2(new_n727), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n987), .B(new_n1147), .C1(new_n418), .C2(new_n731), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n735), .A2(new_n251), .B1(new_n738), .B2(new_n758), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n747), .A2(new_n205), .B1(new_n744), .B2(new_n559), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1148), .A2(new_n946), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT58), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT58), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1146), .B(new_n362), .C1(G33), .C2(G41), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n725), .A2(new_n1063), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n789), .A2(G132), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G128), .A2(new_n727), .B1(new_n730), .B2(G137), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n792), .A2(G125), .B1(new_n793), .B2(G150), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n261), .B(new_n316), .C1(new_n735), .C2(new_n947), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G124), .B2(new_n739), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n715), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n703), .C1(G50), .C2(new_n787), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1127), .B2(new_n712), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n702), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1170), .ZN(G375));
  NAND2_X1  g0971(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1087), .A2(new_n712), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n703), .B1(G68), .B2(new_n787), .ZN(new_n1174));
  INV_X1    g0974(.A(G128), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n731), .A2(new_n801), .B1(new_n738), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G137), .B2(new_n727), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n725), .A2(G159), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n268), .B1(new_n735), .B2(new_n251), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n789), .B2(new_n1063), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n792), .A2(G132), .B1(new_n793), .B2(G50), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n731), .A2(new_n206), .B1(new_n761), .B2(new_n744), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G116), .B2(new_n789), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT123), .Z(new_n1185));
  NAND2_X1  g0985(.A1(new_n950), .A2(new_n265), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT124), .Z(new_n1187));
  NOR2_X1   g0987(.A1(new_n738), .A2(new_n570), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1188), .B(new_n988), .C1(G283), .C2(new_n727), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n205), .C2(new_n724), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1182), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1174), .B1(new_n1191), .B2(new_n715), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1172), .A2(new_n702), .B1(new_n1173), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1107), .A2(new_n927), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1104), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G381));
  INV_X1    g0998(.A(G375), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1015), .A2(new_n769), .A3(new_n1016), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n784), .A2(new_n814), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1050), .A2(new_n1201), .A3(new_n1197), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(G387), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G378), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1199), .A2(new_n1203), .A3(new_n1204), .ZN(G407));
  NAND3_X1  g1005(.A1(new_n620), .A2(new_n621), .A3(G213), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1199), .A2(new_n1204), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(G407), .A2(new_n1208), .A3(G213), .ZN(G409));
  NAND2_X1  g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1200), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n945), .A2(new_n971), .A3(G390), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G390), .B1(new_n945), .B2(new_n971), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1211), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1145), .A2(G378), .A3(new_n1170), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1170), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1139), .A2(new_n927), .A3(new_n1141), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1099), .B1(new_n1116), .B2(new_n1117), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1107), .A2(new_n1048), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1196), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(KEYINPUT125), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT60), .B1(new_n1196), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G384), .A2(new_n1193), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1193), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1201), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1224), .A2(new_n1225), .A3(new_n1206), .A4(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1207), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1207), .A2(G2897), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1236), .B(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1237), .B(new_n1238), .C1(new_n1239), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1207), .B(new_n1243), .C1(new_n1220), .C2(new_n1223), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(new_n1225), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1219), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1215), .A2(new_n1218), .A3(new_n1238), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1244), .B2(KEYINPUT63), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1224), .A2(new_n1206), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1243), .B(new_n1240), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT126), .B1(new_n1241), .B2(new_n1239), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1249), .B2(new_n1243), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1248), .A2(new_n1252), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1246), .A2(new_n1256), .ZN(G405));
  NAND2_X1  g1057(.A1(G375), .A2(new_n1204), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1220), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1236), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1220), .A3(new_n1243), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1215), .A2(new_n1218), .A3(KEYINPUT127), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT127), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1263), .B(new_n1264), .ZN(G402));
endmodule


