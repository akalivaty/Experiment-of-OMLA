//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(new_n462), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT66), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(KEYINPUT66), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n477), .B2(G101), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n468), .B(new_n473), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(G2105), .A3(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n462), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(G136), .B2(new_n491), .ZN(G162));
  OR2_X1    g067(.A1(new_n472), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n487), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n486), .A2(new_n462), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n486), .A2(new_n503), .A3(new_n462), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  NOR4_X1   g080(.A1(new_n465), .A2(KEYINPUT4), .A3(new_n499), .A4(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n498), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n511), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G166));
  XNOR2_X1  g102(.A(new_n521), .B(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n530), .B2(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n531), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n521), .B(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  INV_X1    g118(.A(new_n522), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT71), .B(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(new_n545), .B1(G52), .B2(new_n515), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n511), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n515), .A2(G43), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT72), .B(G81), .Z(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n522), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n515), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n521), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G651), .A2(new_n566), .B1(new_n544), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G166), .ZN(G303));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n511), .B1(new_n540), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G49), .B2(new_n515), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n544), .A2(G87), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G288));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n519), .B2(new_n520), .ZN(new_n578));
  AND2_X1   g153(.A1(G73), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n515), .A2(G48), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(G86), .A3(new_n521), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT75), .Z(G305));
  AOI22_X1  g159(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n511), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n515), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n522), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  NAND3_X1  g167(.A1(G301), .A2(new_n592), .A3(G868), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n564), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT10), .B1(new_n544), .B2(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n592), .B1(G301), .B2(G868), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n594), .B1(new_n603), .B2(new_n604), .ZN(G284));
  AOI21_X1  g180(.A(new_n594), .B1(new_n603), .B2(new_n604), .ZN(G321));
  NOR2_X1   g181(.A1(G286), .A2(new_n602), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n562), .A2(new_n567), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT77), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n602), .ZN(G297));
  AOI21_X1  g185(.A(new_n607), .B1(new_n609), .B2(new_n602), .ZN(G280));
  INV_X1    g186(.A(new_n601), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(new_n465), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n477), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n491), .A2(G135), .ZN(new_n624));
  INV_X1    g199(.A(new_n487), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n472), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n624), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT78), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n622), .A2(G2100), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n623), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT79), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n638), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n646), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT80), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n653), .B(new_n654), .C1(new_n442), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(KEYINPUT81), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n442), .A2(new_n655), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n653), .A2(new_n658), .A3(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  AOI211_X1 g251(.A(new_n674), .B(new_n676), .C1(new_n669), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(G1981), .B(G1986), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G33), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT25), .Z(new_n688));
  AOI22_X1  g263(.A1(new_n619), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n689));
  INV_X1    g264(.A(G139), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n471), .A2(new_n472), .ZN(new_n691));
  OAI221_X1 g266(.A(new_n688), .B1(new_n689), .B2(new_n472), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT90), .Z(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n686), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2072), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT24), .B(G34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(new_n694), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n482), .B2(new_n694), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT27), .B(G1996), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n491), .A2(G141), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT26), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n477), .A2(G105), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n708), .B(new_n709), .C1(new_n625), .C2(G129), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n712), .B(new_n713), .C1(G29), .C2(G32), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n696), .B1(new_n697), .B2(new_n701), .C1(new_n703), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n694), .A2(G27), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G164), .B2(new_n694), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G2078), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n722), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G1966), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(G1966), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n694), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n629), .B2(new_n694), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n725), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n722), .A2(G20), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT23), .Z(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT97), .B(G1956), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n491), .A2(G140), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n625), .A2(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n472), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n694), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT88), .B(G2067), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G171), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT95), .B(G1961), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n732), .A2(new_n737), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT86), .Z(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n601), .B2(new_n722), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT87), .B(G1348), .Z(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT29), .B(G2090), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n758), .B(new_n759), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n722), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n554), .B2(new_n722), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n765), .A2(G1341), .B1(new_n761), .B2(new_n762), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n701), .A2(new_n697), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(G1341), .C2(new_n765), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n753), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n715), .A2(new_n703), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  INV_X1    g346(.A(new_n720), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n717), .A2(new_n721), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  MUX2_X1   g349(.A(G6), .B(G305), .S(G16), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n722), .A2(G23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G288), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT33), .B(G1976), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT85), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n722), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n722), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1971), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n779), .B2(new_n781), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n777), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n694), .A2(G25), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n491), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n625), .A2(G119), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n472), .A2(G107), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT84), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n722), .A2(G24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n590), .B2(new_n722), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n798), .A2(new_n799), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n789), .A2(new_n790), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT36), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n774), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(G311));
  XNOR2_X1  g384(.A(new_n808), .B(KEYINPUT98), .ZN(G150));
  NAND2_X1  g385(.A1(new_n528), .A2(G67), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n511), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n515), .A2(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n522), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n813), .A2(KEYINPUT99), .A3(new_n816), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n554), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(KEYINPUT99), .C1(new_n550), .C2(new_n553), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT38), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n612), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  INV_X1    g401(.A(G860), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n813), .A2(new_n816), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(G145));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n625), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n472), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G142), .B2(new_n491), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n621), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n796), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n711), .B(new_n742), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n503), .B1(new_n471), .B2(new_n500), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n507), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n846));
  INV_X1    g421(.A(new_n498), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n842), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n692), .ZN(new_n853));
  INV_X1    g428(.A(new_n851), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n842), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n693), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n841), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G160), .B(new_n629), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G162), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n693), .ZN(new_n861));
  INV_X1    g436(.A(new_n841), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n861), .B(new_n862), .C1(new_n692), .C2(new_n852), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n858), .B2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n834), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n869), .A2(KEYINPUT101), .A3(new_n865), .A4(new_n864), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n608), .A2(new_n601), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT102), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n608), .A2(new_n601), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n875), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n873), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n876), .A2(new_n873), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n822), .B(new_n615), .ZN(new_n885));
  MUX2_X1   g460(.A(new_n882), .B(new_n884), .S(new_n885), .Z(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n590), .B(G305), .ZN(new_n889));
  OR2_X1    g464(.A1(G166), .A2(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(G166), .A2(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(G288), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G288), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT42), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  INV_X1    g476(.A(new_n889), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(KEYINPUT104), .A3(new_n896), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n899), .B1(new_n906), .B2(KEYINPUT42), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n888), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n886), .A2(new_n887), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g488(.A(new_n912), .B1(G868), .B2(new_n830), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n884), .A2(new_n878), .B1(new_n874), .B2(new_n880), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  XNOR2_X1  g492(.A(G286), .B(G301), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n822), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n822), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G286), .B(G171), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n821), .A3(new_n820), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n884), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n822), .A2(new_n918), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n906), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n924), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n922), .A2(new_n926), .B1(new_n882), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n906), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n865), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n915), .B1(new_n934), .B2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(new_n921), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n926), .A2(new_n936), .A3(new_n919), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n882), .A2(new_n930), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n937), .A2(new_n938), .B1(new_n905), .B2(new_n901), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT107), .B1(new_n939), .B2(G37), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n865), .C1(new_n931), .C2(new_n932), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n942), .A3(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n935), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n929), .A2(new_n947), .A3(new_n865), .A4(new_n933), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n945), .B1(new_n949), .B2(new_n915), .ZN(new_n950));
  AOI211_X1 g525(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n946), .C2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n950), .B2(new_n951), .ZN(G397));
  XNOR2_X1  g527(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n851), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G40), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n482), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT110), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n742), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n711), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(new_n963), .A3(new_n711), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n799), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n797), .A2(new_n968), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n967), .A2(new_n969), .B1(G2067), .B2(new_n742), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(new_n960), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n959), .A2(new_n963), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT46), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n962), .A2(new_n711), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n960), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n796), .B(new_n968), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n967), .B1(new_n960), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1986), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n959), .A2(new_n980), .A3(new_n590), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT48), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n971), .B(new_n977), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n845), .B2(new_n847), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n958), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n954), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT117), .B(new_n958), .C1(new_n984), .C2(KEYINPUT45), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n958), .B1(new_n984), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n506), .B1(new_n994), .B2(new_n502), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n992), .B(new_n955), .C1(new_n995), .C2(new_n498), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT112), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n984), .A2(new_n998), .A3(new_n992), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n990), .A2(new_n991), .B1(new_n1000), .B2(new_n697), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT124), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n989), .A2(new_n988), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT117), .B1(new_n1006), .B2(new_n958), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n991), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G160), .A2(G40), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n955), .B1(new_n995), .B2(new_n498), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(KEYINPUT50), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n998), .B1(new_n984), .B2(new_n992), .ZN(new_n1012));
  NOR4_X1   g587(.A1(G164), .A2(KEYINPUT112), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1011), .B(new_n697), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1002), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n1002), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(KEYINPUT51), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1003), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT51), .B(G8), .C1(new_n1021), .C2(G286), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1015), .C2(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(new_n1018), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1030), .A3(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT55), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(new_n953), .C1(G164), .C2(G1384), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n958), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n1010), .B2(new_n953), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT100), .B1(new_n995), .B2(new_n498), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(KEYINPUT45), .A3(new_n955), .A4(new_n848), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1971), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G2090), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1011), .B(new_n1043), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1034), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1002), .B1(new_n984), .B2(new_n958), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n572), .A2(new_n575), .A3(G1976), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n583), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT116), .B1(new_n583), .B2(G1981), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT114), .B(G1981), .Z(new_n1055));
  NAND4_X1  g630(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT115), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1056), .B(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(KEYINPUT49), .C1(new_n1053), .C2(new_n1052), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1061), .A3(new_n1047), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1065), .A2(new_n1047), .A3(KEYINPUT113), .A4(new_n1048), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1043), .A2(new_n1071), .A3(new_n996), .A4(new_n958), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT111), .B1(new_n984), .B2(new_n954), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1041), .A2(new_n958), .A3(new_n1073), .A4(new_n1036), .ZN(new_n1074));
  INV_X1    g649(.A(G1971), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1033), .B1(new_n1076), .B2(new_n1002), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1046), .A2(new_n1070), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1074), .B2(G2078), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(G2078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT125), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1079), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1029), .A2(new_n1031), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  INV_X1    g669(.A(new_n996), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n993), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n562), .A2(new_n1097), .A3(new_n567), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n562), .B2(new_n567), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1096), .B(new_n1101), .C1(new_n1074), .C2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1100), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1098), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1036), .A2(new_n958), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(new_n1041), .A3(new_n1073), .A4(new_n1102), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT120), .B(new_n1109), .C1(new_n1111), .C2(new_n1096), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1096), .B1(new_n1074), .B2(new_n1103), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1109), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n984), .A2(new_n961), .A3(new_n958), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1000), .B2(G1348), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(new_n612), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1104), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT60), .B(new_n1118), .C1(new_n1000), .C2(G1348), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n612), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n601), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1127), .A2(new_n1128), .B1(new_n1129), .B2(new_n1119), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1074), .B2(G1996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n554), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1136), .A3(new_n554), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1104), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1101), .B1(new_n1111), .B2(new_n1096), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1104), .A2(KEYINPUT121), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1111), .A2(new_n1144), .A3(new_n1096), .A4(new_n1101), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1138), .B(new_n1142), .C1(new_n1117), .C2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1121), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1073), .A2(new_n958), .A3(new_n1036), .ZN(new_n1149));
  AND4_X1   g724(.A1(KEYINPUT45), .A2(new_n1040), .A3(new_n955), .A4(new_n848), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT53), .B1(new_n1151), .B2(new_n771), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n468), .A2(G40), .A3(new_n1082), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n478), .B(KEYINPUT67), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n473), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT126), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1157), .A3(new_n473), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1041), .A2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1000), .A2(G1961), .B1(new_n956), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(G171), .B1(new_n1152), .B2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1081), .A2(G301), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(KEYINPUT54), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1078), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n1166));
  OR3_X1    g741(.A1(new_n1152), .A2(new_n1161), .A3(G171), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1089), .A2(new_n1091), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1148), .A2(new_n1169), .A3(new_n1028), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1062), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(G1976), .A3(G288), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1047), .B1(new_n1172), .B2(new_n1057), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1070), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1046), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1001), .A2(new_n1002), .A3(G286), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1176), .A2(KEYINPUT63), .A3(new_n1046), .ZN(new_n1177));
  OAI21_X1  g752(.A(G8), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1033), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(new_n1070), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1180), .B1(new_n1179), .B2(new_n1070), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1177), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1078), .A2(new_n1176), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1175), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1093), .A2(new_n1170), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n590), .B(new_n980), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n959), .A2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n979), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1190), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n983), .B1(new_n1194), .B2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(G319), .ZN(new_n1198));
  NOR4_X1   g772(.A1(G229), .A2(new_n1198), .A3(G401), .A4(G227), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n871), .A2(new_n949), .A3(new_n1199), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


