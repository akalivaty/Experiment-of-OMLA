//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT86), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT86), .A2(G143), .ZN(new_n190));
  OAI211_X1 g004(.A(G214), .B(new_n188), .C1(new_n189), .C2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G214), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT86), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n198), .A2(new_n199), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n200), .A3(new_n202), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT74), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G140), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(new_n210), .B2(G125), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT74), .A3(G125), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G125), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G140), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n213), .B2(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT89), .B1(new_n206), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n202), .B1(new_n197), .B2(new_n200), .ZN(new_n225));
  AOI211_X1 g039(.A(new_n199), .B(new_n198), .C1(new_n191), .C2(new_n196), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n213), .A2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT88), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n220), .A3(new_n215), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT16), .B1(new_n210), .B2(G125), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n219), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI211_X1 g051(.A(G146), .B(new_n235), .C1(new_n213), .C2(KEYINPUT16), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n191), .B2(new_n196), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT17), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n197), .A2(G131), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n243), .A2(new_n241), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n239), .B(new_n242), .C1(new_n244), .C2(KEYINPUT17), .ZN(new_n245));
  XNOR2_X1  g059(.A(G113), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(G104), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n233), .B2(new_n245), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n187), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G475), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G122), .ZN(new_n261));
  INV_X1    g075(.A(G107), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G116), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT14), .A3(G122), .ZN(new_n265));
  INV_X1    g079(.A(new_n261), .ZN(new_n266));
  OAI211_X1 g080(.A(G107), .B(new_n265), .C1(new_n266), .C2(KEYINPUT14), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n255), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n257), .B1(new_n269), .B2(KEYINPUT13), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n255), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G134), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n261), .B(new_n262), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n259), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT9), .B(G234), .ZN(new_n278));
  INV_X1    g092(.A(G217), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n278), .A2(new_n279), .A3(G953), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n268), .A2(new_n276), .A3(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G478), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT15), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n187), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n193), .A2(G952), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(G237), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n187), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT21), .B(G898), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n287), .B1(new_n284), .B2(new_n187), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n235), .B1(new_n213), .B2(KEYINPUT16), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n243), .A2(new_n241), .B1(new_n298), .B2(new_n219), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n213), .A2(KEYINPUT19), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n216), .A2(new_n218), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(KEYINPUT19), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G146), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n224), .B2(new_n232), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n297), .B1(new_n305), .B2(new_n248), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n299), .A2(new_n303), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n228), .B1(new_n227), .B2(new_n231), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n248), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(KEYINPUT90), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n312), .A3(new_n249), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n314));
  NOR2_X1   g128(.A1(G475), .A2(G902), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n253), .B(new_n296), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT20), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(KEYINPUT91), .A3(new_n253), .A4(new_n296), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G469), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT12), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT11), .B1(new_n259), .B2(G137), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT11), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n333), .B2(G134), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n259), .A2(KEYINPUT65), .A3(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n335), .A2(new_n240), .A3(new_n337), .A4(new_n338), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n219), .A2(G143), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n254), .A2(G146), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n219), .A2(KEYINPUT64), .A3(G143), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT64), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n254), .B2(G146), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n254), .A2(G146), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(KEYINPUT1), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G128), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n345), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n262), .A3(G104), .ZN(new_n356));
  INV_X1    g170(.A(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n247), .A2(G107), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n247), .A2(G107), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n262), .A2(G104), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n351), .A2(G128), .B1(new_n343), .B2(new_n344), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n359), .B(new_n362), .C1(new_n365), .C2(new_n345), .ZN(new_n366));
  AOI221_X4 g180(.A(new_n330), .B1(new_n340), .B2(new_n341), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n340), .A2(new_n341), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT12), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n350), .A2(new_n352), .ZN(new_n372));
  INV_X1    g186(.A(new_n345), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n359), .A2(new_n362), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT10), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT0), .A2(G128), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n343), .A2(new_n344), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n350), .A2(new_n384), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n387), .A3(G101), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n341), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n337), .A2(new_n338), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n240), .B1(new_n391), .B2(new_n335), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n376), .A2(new_n378), .A3(new_n389), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n193), .A2(G227), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT80), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G140), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n371), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n376), .A2(new_n378), .A3(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n369), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n398), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n329), .B(new_n187), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n329), .A2(new_n187), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n394), .B1(new_n367), .B2(new_n370), .ZN(new_n407));
  INV_X1    g221(.A(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n394), .A2(new_n398), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n402), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(G469), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n404), .A2(new_n406), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G221), .B1(new_n278), .B2(G902), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT79), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(G224), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n384), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n344), .A2(KEYINPUT64), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n343), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n424), .B2(new_n346), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n385), .A2(new_n382), .ZN(new_n426));
  OAI21_X1  g240(.A(G125), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n353), .A2(new_n217), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n427), .A2(new_n419), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n375), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n264), .A2(G119), .ZN(new_n435));
  INV_X1    g249(.A(G119), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT67), .B1(new_n436), .B2(G116), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n264), .A3(G119), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT2), .B(G113), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n439), .ZN(new_n443));
  INV_X1    g257(.A(new_n435), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(KEYINPUT5), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G113), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n434), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT8), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n442), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(KEYINPUT85), .B2(new_n363), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n450), .B(new_n452), .C1(new_n454), .C2(new_n434), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n427), .A2(new_n428), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n420), .A3(new_n419), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n431), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n375), .A3(new_n442), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n440), .A2(new_n441), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n388), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n451), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n440), .B(new_n441), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n381), .A3(new_n388), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n451), .A4(new_n459), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n187), .B1(new_n458), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n469), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n451), .B1(new_n467), .B2(new_n459), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n429), .A2(new_n430), .ZN(new_n479));
  AOI211_X1 g293(.A(KEYINPUT6), .B(new_n451), .C1(new_n467), .C2(new_n459), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n473), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n474), .B2(new_n477), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n473), .B1(new_n483), .B2(new_n479), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n481), .A3(new_n479), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n473), .A3(new_n479), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n486), .A3(new_n472), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n328), .B(new_n417), .C1(new_n488), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n188), .A2(G210), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT27), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n333), .B2(G134), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n333), .A2(G134), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n259), .A2(KEYINPUT66), .A3(G137), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G131), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n341), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n341), .A2(KEYINPUT68), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n374), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n466), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT28), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n353), .B1(new_n506), .B2(new_n507), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n515), .A2(new_n509), .B1(new_n369), .B2(new_n386), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n374), .A2(new_n341), .A3(new_n505), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n512), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n466), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n499), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n510), .B2(new_n512), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n512), .A3(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n466), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n513), .A3(new_n499), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n528), .A2(KEYINPUT31), .A3(new_n513), .A4(new_n499), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT32), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n495), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT69), .B(KEYINPUT32), .Z(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n533), .B2(new_n535), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n519), .A2(new_n522), .A3(new_n499), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  INV_X1    g357(.A(new_n513), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n526), .B1(new_n516), .B2(new_n524), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n466), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n542), .B(new_n543), .C1(new_n546), .C2(new_n499), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n516), .A2(new_n511), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n514), .B2(new_n518), .ZN(new_n549));
  INV_X1    g363(.A(new_n499), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n543), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  INV_X1    g368(.A(new_n523), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT31), .B1(new_n546), .B2(new_n499), .ZN(new_n556));
  AND4_X1   g370(.A1(KEYINPUT31), .A2(new_n528), .A3(new_n513), .A4(new_n499), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT70), .A3(new_n537), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n539), .A2(new_n541), .A3(new_n554), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT76), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT22), .B(G137), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n436), .B2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n436), .A2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n256), .A2(KEYINPUT71), .A3(G119), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT24), .B(G110), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n436), .B2(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT72), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n575), .A2(new_n576), .A3(new_n579), .A4(new_n568), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n573), .A2(new_n578), .A3(G110), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G110), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n577), .B2(KEYINPUT72), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n573), .B1(new_n583), .B2(new_n580), .ZN(new_n584));
  OAI221_X1 g398(.A(new_n572), .B1(new_n237), .B2(new_n238), .C1(new_n581), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n571), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(G110), .B2(new_n577), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n587), .B(new_n220), .C1(new_n219), .C2(new_n298), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n565), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n581), .A2(new_n584), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n572), .B1(new_n237), .B2(new_n238), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n565), .B(new_n588), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n564), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n564), .B1(new_n595), .B2(KEYINPUT77), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n187), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT78), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT25), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n592), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n596), .B1(new_n603), .B2(new_n564), .ZN(new_n604));
  INV_X1    g418(.A(new_n600), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n187), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n279), .B1(G234), .B2(new_n187), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(G902), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n607), .A2(new_n608), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n326), .A2(new_n494), .A3(new_n560), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  OAI21_X1  g426(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n558), .A2(new_n534), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n605), .B1(new_n604), .B2(new_n187), .ZN(new_n616));
  INV_X1    g430(.A(new_n564), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n602), .B2(new_n592), .ZN(new_n618));
  NOR4_X1   g432(.A1(new_n618), .A2(G902), .A3(new_n596), .A4(new_n600), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n608), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n604), .A2(new_n609), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n615), .A2(new_n622), .A3(new_n417), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT92), .Z(new_n624));
  AOI21_X1  g438(.A(new_n328), .B1(new_n488), .B2(new_n493), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n253), .B1(new_n316), .B2(new_n317), .ZN(new_n626));
  INV_X1    g440(.A(new_n294), .ZN(new_n627));
  INV_X1    g441(.A(new_n283), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n280), .B1(new_n268), .B2(new_n276), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n285), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n285), .A2(new_n187), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n628), .B2(KEYINPUT93), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n630), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n632), .B(new_n634), .C1(new_n636), .C2(new_n285), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n624), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NOR2_X1   g457(.A1(new_n289), .A2(new_n295), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n252), .B2(G475), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n294), .B(KEYINPUT94), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n625), .A2(new_n324), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n624), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT95), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n595), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n609), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n607), .B2(new_n608), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT96), .B1(new_n615), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n620), .A2(new_n655), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n614), .A4(new_n613), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n326), .A2(new_n658), .A3(new_n494), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G12));
  XOR2_X1   g479(.A(new_n291), .B(KEYINPUT98), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n292), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n645), .B(new_n670), .C1(new_n316), .C2(new_n317), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n494), .A2(new_n560), .A3(new_n659), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  AND2_X1   g488(.A1(new_n539), .A2(new_n559), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n546), .A2(new_n550), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n513), .A2(new_n550), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n187), .B1(new_n677), .B2(new_n548), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n675), .A2(new_n541), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n488), .A2(new_n493), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n682), .B1(new_n488), .B2(new_n493), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n669), .B(KEYINPUT39), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n417), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n407), .A2(new_n408), .B1(new_n410), .B2(new_n402), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n405), .B1(new_n690), .B2(G469), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n415), .B1(new_n691), .B2(new_n404), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT100), .B1(new_n692), .B2(new_n687), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  OAI221_X1 g509(.A(new_n680), .B1(new_n684), .B2(new_n685), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n644), .B1(new_n324), .B2(new_n253), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(new_n327), .A3(new_n657), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n254), .ZN(G45));
  AOI22_X1  g515(.A1(new_n614), .A2(new_n540), .B1(G472), .B2(new_n553), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n657), .B1(new_n675), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n626), .A2(new_n638), .A3(new_n670), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n626), .A2(new_n638), .A3(KEYINPUT101), .A4(new_n670), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n494), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  OAI21_X1  g523(.A(new_n187), .B1(new_n400), .B2(new_n403), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n416), .A3(new_n404), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n560), .A2(new_n610), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n639), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT102), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n715), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n714), .A2(new_n647), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n264), .ZN(G18));
  AOI211_X1 g534(.A(new_n328), .B(new_n712), .C1(new_n488), .C2(new_n493), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n326), .A2(new_n721), .A3(new_n560), .A4(new_n659), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n703), .A2(new_n724), .A3(new_n326), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  INV_X1    g541(.A(new_n548), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n499), .B1(new_n519), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n531), .B2(new_n532), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT104), .B1(new_n730), .B2(new_n535), .ZN(new_n731));
  INV_X1    g545(.A(new_n729), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n556), .B2(new_n557), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n534), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n613), .A2(KEYINPUT105), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(G472), .C1(new_n533), .C2(G902), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n737), .A3(new_n610), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n625), .A2(new_n713), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n698), .A2(new_n646), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(G122), .Z(G24));
  AND4_X1   g558(.A1(new_n659), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n706), .A3(new_n707), .A4(new_n721), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT106), .B(G125), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G27));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n706), .A2(new_n707), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n488), .A2(new_n493), .A3(new_n327), .A4(new_n692), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n560), .A3(new_n610), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n749), .ZN(new_n755));
  AOI22_X1  g569(.A1(G472), .A2(new_n553), .B1(new_n558), .B2(new_n537), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n614), .A2(new_n536), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n622), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n706), .A3(new_n758), .A4(new_n707), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n671), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n671), .B(KEYINPUT107), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n622), .B1(new_n675), .B2(new_n702), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT108), .A4(new_n752), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NOR2_X1   g584(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n329), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n405), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n404), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT109), .A3(new_n416), .A4(new_n687), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n416), .B1(new_n775), .B2(new_n776), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n779), .B1(new_n780), .B2(new_n688), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n488), .A2(new_n493), .A3(new_n327), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n778), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n615), .A2(new_n659), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT110), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n324), .A2(new_n253), .A3(new_n638), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n786), .A2(new_n791), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n784), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT111), .B(G137), .Z(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n780), .B(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n706), .A2(new_n707), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n560), .A2(new_n782), .A3(new_n610), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n711), .A2(new_n404), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n328), .B(new_n415), .C1(new_n805), .C2(KEYINPUT49), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(KEYINPUT49), .B2(new_n805), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n622), .A3(new_n787), .ZN(new_n808));
  INV_X1    g622(.A(new_n680), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n684), .A2(new_n685), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n714), .B1(new_n639), .B2(new_n647), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n743), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n726), .ZN(new_n814));
  INV_X1    g628(.A(new_n646), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n328), .B(new_n815), .C1(new_n488), .C2(new_n493), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n626), .A2(new_n638), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n324), .A2(new_n645), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n623), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n662), .A2(new_n611), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n662), .A2(new_n611), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n324), .A2(new_n253), .A3(new_n644), .A4(new_n670), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n751), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n703), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n706), .A2(new_n707), .A3(new_n752), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n736), .A2(new_n737), .A3(new_n659), .A4(new_n739), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n754), .B2(new_n759), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n814), .A2(new_n825), .A3(new_n769), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n486), .B1(new_n492), .B2(new_n472), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n487), .B(new_n471), .C1(new_n490), .C2(new_n491), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n327), .B(new_n692), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n626), .B1(new_n295), .B2(new_n289), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n620), .A2(new_n655), .A3(new_n670), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT114), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n620), .A2(new_n841), .A3(new_n655), .A4(new_n670), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n838), .A2(new_n843), .A3(new_n680), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n746), .A2(new_n708), .A3(new_n673), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n494), .A2(new_n560), .A3(new_n659), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n801), .B2(new_n672), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n746), .A4(new_n844), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n833), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n855), .B(new_n854), .C1(new_n833), .C2(new_n851), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n290), .B(KEYINPUT118), .Z(new_n861));
  NOR2_X1   g675(.A1(new_n782), .A2(new_n712), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n610), .A2(new_n291), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n809), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n864), .B2(new_n817), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n740), .A2(new_n741), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n666), .B1(new_n789), .B2(new_n790), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n758), .A3(new_n862), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT48), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT48), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n871), .A3(new_n758), .A4(new_n862), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n868), .A2(new_n873), .A3(KEYINPUT119), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT119), .B1(new_n868), .B2(new_n873), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n740), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n712), .A2(new_n327), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n867), .A2(new_n877), .A3(new_n810), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n324), .A2(new_n253), .A3(new_n637), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n809), .A2(new_n862), .A3(new_n863), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n867), .A2(new_n862), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n830), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n867), .A2(new_n877), .A3(new_n783), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n780), .B(KEYINPUT47), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n805), .A2(new_n416), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT116), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n889), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n884), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n899));
  OAI211_X1 g713(.A(KEYINPUT51), .B(new_n887), .C1(new_n888), .C2(new_n830), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n890), .B1(new_n800), .B2(new_n892), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n882), .A3(new_n883), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n876), .A2(new_n898), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n855), .B1(new_n833), .B2(new_n851), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT115), .B1(new_n813), .B2(new_n726), .ZN(new_n906));
  INV_X1    g720(.A(new_n829), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n907), .A2(new_n745), .B1(new_n703), .B2(new_n827), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n760), .A2(new_n908), .A3(new_n769), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n846), .A2(new_n850), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n855), .B1(new_n822), .B2(new_n824), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n905), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n903), .B1(new_n874), .B2(new_n875), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT51), .B1(new_n884), .B2(new_n895), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT120), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n860), .A2(new_n904), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n811), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n193), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n187), .B1(new_n905), .B2(new_n914), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n483), .B(new_n479), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n926), .B2(new_n929), .ZN(G51));
  INV_X1    g745(.A(new_n916), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n915), .B1(new_n905), .B2(new_n914), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n405), .B(KEYINPUT57), .Z(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n403), .B2(new_n400), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n773), .A3(new_n772), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n923), .B1(new_n936), .B2(new_n937), .ZN(G54));
  AND3_X1   g752(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(new_n313), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n924), .B1(new_n939), .B2(new_n313), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(new_n860), .A2(new_n916), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n633), .B(KEYINPUT59), .Z(new_n944));
  AOI21_X1  g758(.A(new_n636), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n636), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n924), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(new_n905), .A2(new_n914), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT121), .Z(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n604), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n923), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  INV_X1    g771(.A(new_n952), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n905), .B2(new_n914), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n654), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n956), .A2(new_n957), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n924), .B1(new_n959), .B2(new_n604), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n949), .A2(new_n654), .A3(new_n952), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n962), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n961), .A2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n293), .B2(new_n418), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n814), .A2(new_n825), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n970), .B2(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n483), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(G898), .B2(new_n193), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n625), .A2(new_n698), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n778), .A2(new_n781), .A3(new_n758), .A4(new_n977), .ZN(new_n978));
  AND4_X1   g792(.A1(new_n760), .A2(new_n803), .A3(new_n769), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n494), .A2(new_n560), .A3(new_n659), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n673), .B1(new_n980), .B2(new_n750), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n750), .A2(new_n741), .A3(new_n830), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT123), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n746), .A2(new_n708), .A3(new_n984), .A4(new_n673), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n979), .A2(new_n193), .A3(new_n796), .A4(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n545), .B(new_n302), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(G900), .B2(G953), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n987), .A2(new_n989), .B1(KEYINPUT126), .B2(new_n975), .ZN(new_n990));
  INV_X1    g804(.A(new_n988), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n767), .A2(new_n694), .A3(new_n783), .A4(new_n819), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n801), .A2(new_n802), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n994), .B(new_n995), .C1(new_n891), .C2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n778), .A2(new_n781), .A3(new_n783), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n794), .B2(new_n793), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n997), .B1(new_n999), .B2(new_n792), .ZN(new_n1000));
  INV_X1    g814(.A(new_n700), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT62), .B1(new_n986), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n1003), .B(new_n700), .C1(new_n983), .C2(new_n985), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n991), .B1(new_n1005), .B2(new_n193), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT125), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n990), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g822(.A(KEYINPUT125), .B(new_n991), .C1(new_n1005), .C2(new_n193), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n976), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n796), .A2(new_n803), .A3(new_n994), .A4(new_n995), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n986), .A2(new_n1001), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n1003), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n986), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n988), .B1(new_n1015), .B2(G953), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .ZN(new_n1017));
  INV_X1    g831(.A(new_n976), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n990), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1010), .A2(new_n1020), .ZN(G72));
  INV_X1    g835(.A(new_n528), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n677), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND3_X1  g839(.A1(new_n979), .A2(new_n796), .A3(new_n986), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n969), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1027), .A2(KEYINPUT127), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1029), .B(new_n1025), .C1(new_n1026), .C2(new_n969), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1023), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1015), .A2(new_n970), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1025), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n676), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n550), .B1(new_n1022), .B2(new_n544), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1035), .B1(new_n1037), .B2(new_n529), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n923), .B1(new_n859), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1032), .A2(new_n1036), .A3(new_n1039), .ZN(G57));
endmodule


