

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805;

  NAND2_X2 U375 ( .A1(n539), .A2(n538), .ZN(n541) );
  XNOR2_X2 U376 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X2 U377 ( .A(n738), .B(n737), .ZN(n739) );
  OR2_X2 U378 ( .A1(n746), .A2(G902), .ZN(n466) );
  NOR2_X2 U379 ( .A1(n706), .A2(n716), .ZN(n422) );
  NAND2_X1 U380 ( .A1(n608), .A2(n594), .ZN(n595) );
  XNOR2_X1 U381 ( .A(n388), .B(KEYINPUT30), .ZN(n608) );
  NAND2_X2 U382 ( .A1(n357), .A2(n356), .ZN(n395) );
  INV_X1 U383 ( .A(n452), .ZN(n356) );
  INV_X1 U384 ( .A(n619), .ZN(n357) );
  NOR2_X1 U385 ( .A1(n804), .A2(n557), .ZN(n558) );
  OR2_X2 U386 ( .A1(n535), .A2(n614), .ZN(n672) );
  AND2_X2 U387 ( .A1(n531), .A2(n530), .ZN(n539) );
  XNOR2_X2 U388 ( .A(n358), .B(n446), .ZN(n619) );
  NOR2_X1 U389 ( .A1(n767), .A2(n758), .ZN(n387) );
  NOR2_X1 U390 ( .A1(n751), .A2(n441), .ZN(n383) );
  BUF_X1 U391 ( .A(n392), .Z(n744) );
  NOR2_X1 U392 ( .A1(n556), .A2(n673), .ZN(n557) );
  NAND2_X1 U393 ( .A1(n389), .A2(n397), .ZN(n551) );
  XNOR2_X1 U394 ( .A(n591), .B(n593), .ZN(n675) );
  XNOR2_X1 U395 ( .A(n383), .B(n384), .ZN(n590) );
  NOR2_X1 U396 ( .A1(n451), .A2(n585), .ZN(n452) );
  XNOR2_X1 U397 ( .A(n445), .B(n444), .ZN(n678) );
  NAND2_X1 U398 ( .A1(n590), .A2(n678), .ZN(n358) );
  BUF_X1 U399 ( .A(n500), .Z(n359) );
  NAND2_X1 U400 ( .A1(n418), .A2(n423), .ZN(n360) );
  NAND2_X1 U401 ( .A1(n418), .A2(n423), .ZN(n417) );
  NOR2_X1 U402 ( .A1(n619), .A2(n452), .ZN(n361) );
  NAND2_X1 U403 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U404 ( .A(n575), .B(n574), .ZN(n580) );
  XNOR2_X1 U405 ( .A(n581), .B(KEYINPUT45), .ZN(n362) );
  XNOR2_X1 U406 ( .A(n581), .B(KEYINPUT45), .ZN(n713) );
  NAND2_X1 U407 ( .A1(n377), .A2(n554), .ZN(n676) );
  INV_X1 U408 ( .A(n555), .ZN(n377) );
  XNOR2_X1 U409 ( .A(n378), .B(G146), .ZN(n473) );
  INV_X1 U410 ( .A(G125), .ZN(n378) );
  XNOR2_X1 U411 ( .A(n413), .B(n412), .ZN(n492) );
  XNOR2_X1 U412 ( .A(G116), .B(G113), .ZN(n412) );
  XNOR2_X1 U413 ( .A(n429), .B(n414), .ZN(n413) );
  INV_X1 U414 ( .A(KEYINPUT71), .ZN(n414) );
  NAND2_X1 U415 ( .A1(n416), .A2(n716), .ZN(n415) );
  XNOR2_X1 U416 ( .A(n400), .B(KEYINPUT41), .ZN(n693) );
  NAND2_X1 U417 ( .A1(n404), .A2(n365), .ZN(n629) );
  XNOR2_X1 U418 ( .A(n615), .B(n405), .ZN(n404) );
  INV_X1 U419 ( .A(KEYINPUT107), .ZN(n405) );
  INV_X1 U420 ( .A(KEYINPUT97), .ZN(n386) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n512) );
  XNOR2_X1 U422 ( .A(n434), .B(KEYINPUT17), .ZN(n435) );
  XNOR2_X1 U423 ( .A(n626), .B(n625), .ZN(n636) );
  INV_X1 U424 ( .A(G237), .ZN(n442) );
  XNOR2_X1 U425 ( .A(n363), .B(n473), .ZN(n789) );
  XNOR2_X1 U426 ( .A(G143), .B(G131), .ZN(n517) );
  XNOR2_X1 U427 ( .A(KEYINPUT67), .B(G101), .ZN(n488) );
  XNOR2_X1 U428 ( .A(G134), .B(G131), .ZN(n458) );
  NOR2_X1 U429 ( .A1(n671), .A2(n376), .ZN(n684) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n447) );
  INV_X1 U431 ( .A(KEYINPUT28), .ZN(n399) );
  INV_X1 U432 ( .A(n676), .ZN(n598) );
  INV_X1 U433 ( .A(KEYINPUT0), .ZN(n396) );
  XNOR2_X1 U434 ( .A(n492), .B(n430), .ZN(n779) );
  XNOR2_X1 U435 ( .A(G107), .B(G104), .ZN(n432) );
  XNOR2_X1 U436 ( .A(KEYINPUT78), .B(G110), .ZN(n431) );
  XNOR2_X1 U437 ( .A(G122), .B(G107), .ZN(n503) );
  XOR2_X1 U438 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n504) );
  XNOR2_X1 U439 ( .A(G134), .B(G116), .ZN(n506) );
  XNOR2_X1 U440 ( .A(n511), .B(n510), .ZN(n555) );
  NOR2_X1 U441 ( .A1(n795), .A2(G952), .ZN(n754) );
  NAND2_X1 U442 ( .A1(n392), .A2(G210), .ZN(n374) );
  INV_X1 U443 ( .A(n754), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n409), .B(n408), .ZN(n802) );
  INV_X1 U445 ( .A(KEYINPUT42), .ZN(n408) );
  NAND2_X1 U446 ( .A1(n618), .A2(n657), .ZN(n772) );
  NOR2_X1 U447 ( .A1(n629), .A2(n403), .ZN(n617) );
  XOR2_X1 U448 ( .A(KEYINPUT10), .B(G140), .Z(n363) );
  XOR2_X1 U449 ( .A(n605), .B(n604), .Z(n364) );
  INV_X1 U450 ( .A(n591), .ZN(n403) );
  AND2_X1 U451 ( .A1(n596), .A2(n678), .ZN(n365) );
  NOR2_X1 U452 ( .A1(n623), .A2(n402), .ZN(n366) );
  AND2_X1 U453 ( .A1(n598), .A2(n678), .ZN(n367) );
  AND2_X1 U454 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n368) );
  XOR2_X1 U455 ( .A(n753), .B(n752), .Z(n369) );
  XNOR2_X1 U456 ( .A(n755), .B(KEYINPUT89), .ZN(n370) );
  XNOR2_X1 U457 ( .A(n371), .B(n370), .ZN(G51) );
  NAND2_X1 U458 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U459 ( .A(n374), .B(n369), .ZN(n373) );
  NAND2_X1 U460 ( .A1(n411), .A2(n769), .ZN(n725) );
  XNOR2_X2 U461 ( .A(n595), .B(KEYINPUT39), .ZN(n411) );
  NAND2_X1 U462 ( .A1(n375), .A2(n693), .ZN(n409) );
  INV_X1 U463 ( .A(n620), .ZN(n375) );
  INV_X1 U464 ( .A(n693), .ZN(n376) );
  INV_X1 U465 ( .A(n554), .ZN(n543) );
  INV_X1 U466 ( .A(n789), .ZN(n515) );
  XNOR2_X1 U467 ( .A(n516), .B(n789), .ZN(n524) );
  BUF_X1 U468 ( .A(n492), .Z(n379) );
  XNOR2_X1 U469 ( .A(n566), .B(KEYINPUT106), .ZN(n380) );
  BUF_X1 U470 ( .A(n590), .Z(n591) );
  XNOR2_X1 U471 ( .A(n603), .B(n399), .ZN(n398) );
  NAND2_X2 U472 ( .A1(n395), .A2(n396), .ZN(n389) );
  BUF_X1 U473 ( .A(n727), .Z(n381) );
  XNOR2_X1 U474 ( .A(n410), .B(n597), .ZN(n727) );
  AND2_X2 U475 ( .A1(n571), .A2(n614), .ZN(n382) );
  XNOR2_X2 U476 ( .A(n605), .B(KEYINPUT1), .ZN(n628) );
  NAND2_X1 U477 ( .A1(n398), .A2(n364), .ZN(n620) );
  NAND2_X1 U478 ( .A1(n443), .A2(G210), .ZN(n384) );
  AND2_X1 U479 ( .A1(n394), .A2(n385), .ZN(n758) );
  AND2_X1 U480 ( .A1(n553), .A2(n605), .ZN(n385) );
  XNOR2_X1 U481 ( .A(n387), .B(n386), .ZN(n556) );
  BUF_X1 U482 ( .A(n767), .Z(n770) );
  NOR2_X1 U483 ( .A1(n602), .A2(n599), .ZN(n388) );
  XNOR2_X1 U484 ( .A(n541), .B(n540), .ZN(n576) );
  BUF_X1 U485 ( .A(n459), .Z(n390) );
  BUF_X1 U486 ( .A(n790), .Z(n391) );
  NAND2_X1 U487 ( .A1(n360), .A2(n415), .ZN(n392) );
  NAND2_X1 U488 ( .A1(n397), .A2(n389), .ZN(n393) );
  NAND2_X1 U489 ( .A1(n397), .A2(n389), .ZN(n394) );
  NAND2_X1 U490 ( .A1(n417), .A2(n415), .ZN(n750) );
  NAND2_X1 U491 ( .A1(n361), .A2(KEYINPUT0), .ZN(n397) );
  NAND2_X1 U492 ( .A1(n675), .A2(n598), .ZN(n680) );
  NAND2_X1 U493 ( .A1(n675), .A2(n367), .ZN(n400) );
  NAND2_X1 U494 ( .A1(n772), .A2(n401), .ZN(n402) );
  NOR2_X1 U495 ( .A1(n799), .A2(n368), .ZN(n401) );
  XNOR2_X2 U496 ( .A(n406), .B(G143), .ZN(n500) );
  XNOR2_X2 U497 ( .A(G128), .B(KEYINPUT82), .ZN(n406) );
  XNOR2_X1 U498 ( .A(n407), .B(n493), .ZN(n717) );
  XNOR2_X1 U499 ( .A(n407), .B(n428), .ZN(n746) );
  XNOR2_X2 U500 ( .A(n790), .B(G146), .ZN(n407) );
  NOR2_X2 U501 ( .A1(n727), .A2(n802), .ZN(n606) );
  NAND2_X1 U502 ( .A1(n411), .A2(n596), .ZN(n410) );
  NAND2_X1 U503 ( .A1(n715), .A2(n419), .ZN(n416) );
  NAND2_X1 U504 ( .A1(n421), .A2(n420), .ZN(n418) );
  INV_X1 U505 ( .A(n706), .ZN(n419) );
  INV_X1 U506 ( .A(n424), .ZN(n420) );
  NAND2_X1 U507 ( .A1(n715), .A2(n422), .ZN(n421) );
  NAND2_X1 U508 ( .A1(n424), .A2(KEYINPUT64), .ZN(n423) );
  NOR2_X2 U509 ( .A1(n713), .A2(n702), .ZN(n424) );
  XNOR2_X2 U510 ( .A(n548), .B(n547), .ZN(n571) );
  BUF_X1 U511 ( .A(n576), .Z(n728) );
  XOR2_X1 U512 ( .A(n458), .B(G137), .Z(n425) );
  AND2_X1 U513 ( .A1(n662), .A2(n656), .ZN(n426) );
  AND2_X1 U514 ( .A1(n568), .A2(n659), .ZN(n427) );
  XOR2_X1 U515 ( .A(n462), .B(n461), .Z(n428) );
  XNOR2_X1 U516 ( .A(n435), .B(n473), .ZN(n437) );
  AND2_X1 U517 ( .A1(n582), .A2(n648), .ZN(n653) );
  XNOR2_X1 U518 ( .A(n566), .B(n496), .ZN(n614) );
  BUF_X1 U519 ( .A(n717), .Z(n719) );
  INV_X1 U520 ( .A(KEYINPUT63), .ZN(n723) );
  XNOR2_X1 U521 ( .A(n699), .B(n698), .ZN(G75) );
  INV_X4 U522 ( .A(G953), .ZN(n795) );
  XNOR2_X2 U523 ( .A(G119), .B(KEYINPUT3), .ZN(n429) );
  XNOR2_X1 U524 ( .A(KEYINPUT16), .B(G122), .ZN(n430) );
  XNOR2_X1 U525 ( .A(n432), .B(n431), .ZN(n781) );
  XNOR2_X1 U526 ( .A(n488), .B(KEYINPUT72), .ZN(n433) );
  XNOR2_X1 U527 ( .A(n781), .B(n433), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n779), .B(n462), .ZN(n440) );
  XNOR2_X2 U529 ( .A(n500), .B(KEYINPUT4), .ZN(n459) );
  NAND2_X1 U530 ( .A1(n795), .A2(G224), .ZN(n434) );
  XNOR2_X1 U531 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n436) );
  XNOR2_X1 U532 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U533 ( .A(n390), .B(n438), .ZN(n439) );
  XNOR2_X1 U534 ( .A(n440), .B(n439), .ZN(n751) );
  XNOR2_X1 U535 ( .A(G902), .B(KEYINPUT15), .ZN(n708) );
  INV_X1 U536 ( .A(n708), .ZN(n441) );
  INV_X1 U537 ( .A(G902), .ZN(n525) );
  NAND2_X1 U538 ( .A1(n525), .A2(n442), .ZN(n443) );
  NAND2_X1 U539 ( .A1(n443), .A2(G214), .ZN(n445) );
  INV_X1 U540 ( .A(KEYINPUT93), .ZN(n444) );
  INV_X1 U541 ( .A(KEYINPUT19), .ZN(n446) );
  XNOR2_X1 U542 ( .A(n447), .B(KEYINPUT94), .ZN(n448) );
  XNOR2_X1 U543 ( .A(KEYINPUT14), .B(n448), .ZN(n450) );
  AND2_X1 U544 ( .A1(n450), .A2(G953), .ZN(n449) );
  NAND2_X1 U545 ( .A1(G902), .A2(n449), .ZN(n584) );
  NOR2_X1 U546 ( .A1(n584), .A2(G898), .ZN(n451) );
  NAND2_X1 U547 ( .A1(G952), .A2(n450), .ZN(n688) );
  NOR2_X1 U548 ( .A1(n688), .A2(G953), .ZN(n585) );
  INV_X1 U549 ( .A(KEYINPUT34), .ZN(n498) );
  AND2_X1 U550 ( .A1(n498), .A2(KEYINPUT33), .ZN(n454) );
  NAND2_X1 U551 ( .A1(n551), .A2(n454), .ZN(n457) );
  INV_X1 U552 ( .A(KEYINPUT33), .ZN(n455) );
  NAND2_X1 U553 ( .A1(n455), .A2(KEYINPUT34), .ZN(n456) );
  NAND2_X1 U554 ( .A1(n457), .A2(n456), .ZN(n497) );
  XNOR2_X2 U555 ( .A(n459), .B(n425), .ZN(n790) );
  NAND2_X1 U556 ( .A1(n795), .A2(G227), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n460), .B(G140), .ZN(n461) );
  XNOR2_X1 U558 ( .A(KEYINPUT70), .B(G469), .ZN(n464) );
  INV_X1 U559 ( .A(KEYINPUT69), .ZN(n463) );
  XNOR2_X1 U560 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X2 U561 ( .A(n466), .B(n465), .ZN(n605) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n470) );
  XOR2_X1 U563 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n468) );
  NAND2_X1 U564 ( .A1(G234), .A2(n795), .ZN(n467) );
  XNOR2_X1 U565 ( .A(n468), .B(n467), .ZN(n499) );
  NAND2_X1 U566 ( .A1(G221), .A2(n499), .ZN(n469) );
  XNOR2_X1 U567 ( .A(n470), .B(n469), .ZN(n476) );
  XOR2_X1 U568 ( .A(G110), .B(G119), .Z(n472) );
  XNOR2_X1 U569 ( .A(G128), .B(G137), .ZN(n471) );
  XNOR2_X1 U570 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n474), .B(n515), .ZN(n475) );
  XNOR2_X1 U572 ( .A(n476), .B(n475), .ZN(n729) );
  NAND2_X1 U573 ( .A1(n729), .A2(n525), .ZN(n482) );
  XOR2_X1 U574 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n480) );
  XOR2_X1 U575 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n478) );
  NAND2_X1 U576 ( .A1(G234), .A2(n708), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n483) );
  NAND2_X1 U578 ( .A1(n483), .A2(G217), .ZN(n479) );
  XOR2_X1 U579 ( .A(n480), .B(n479), .Z(n481) );
  XNOR2_X2 U580 ( .A(n482), .B(n481), .ZN(n659) );
  NAND2_X1 U581 ( .A1(G221), .A2(n483), .ZN(n485) );
  INV_X1 U582 ( .A(KEYINPUT21), .ZN(n484) );
  XNOR2_X1 U583 ( .A(n485), .B(n484), .ZN(n660) );
  AND2_X1 U584 ( .A1(n659), .A2(n660), .ZN(n656) );
  NAND2_X1 U585 ( .A1(n628), .A2(n656), .ZN(n535) );
  XOR2_X1 U586 ( .A(KEYINPUT96), .B(KEYINPUT77), .Z(n487) );
  NAND2_X1 U587 ( .A1(n512), .A2(G210), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n488), .B(KEYINPUT5), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n379), .B(n491), .ZN(n493) );
  OR2_X2 U592 ( .A1(n717), .A2(G902), .ZN(n495) );
  XNOR2_X1 U593 ( .A(G472), .B(KEYINPUT73), .ZN(n494) );
  XNOR2_X2 U594 ( .A(n495), .B(n494), .ZN(n566) );
  XNOR2_X1 U595 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n496) );
  NAND2_X1 U596 ( .A1(n497), .A2(n672), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n394), .A2(n498), .ZN(n529) );
  AND2_X1 U598 ( .A1(n499), .A2(G217), .ZN(n502) );
  INV_X1 U599 ( .A(n359), .ZN(n501) );
  XNOR2_X1 U600 ( .A(n502), .B(n501), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U602 ( .A(n505), .B(KEYINPUT101), .Z(n507) );
  XNOR2_X1 U603 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n509), .B(n508), .ZN(n733) );
  NAND2_X1 U605 ( .A1(n733), .A2(n525), .ZN(n511) );
  XNOR2_X1 U606 ( .A(KEYINPUT102), .B(G478), .ZN(n510) );
  XOR2_X1 U607 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n514) );
  NAND2_X1 U608 ( .A1(G214), .A2(n512), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U610 ( .A(G122), .B(G113), .Z(n518) );
  XNOR2_X1 U611 ( .A(n518), .B(n517), .ZN(n522) );
  XOR2_X1 U612 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n520) );
  XNOR2_X1 U613 ( .A(G104), .B(KEYINPUT12), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U616 ( .A(n524), .B(n523), .ZN(n738) );
  NAND2_X1 U617 ( .A1(n738), .A2(n525), .ZN(n527) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  XNOR2_X1 U619 ( .A(n527), .B(n526), .ZN(n554) );
  AND2_X1 U620 ( .A1(n555), .A2(n543), .ZN(n609) );
  INV_X1 U621 ( .A(n609), .ZN(n528) );
  NOR2_X1 U622 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U623 ( .A1(KEYINPUT34), .A2(KEYINPUT33), .ZN(n532) );
  NAND2_X1 U624 ( .A1(n393), .A2(n532), .ZN(n534) );
  NAND2_X1 U625 ( .A1(KEYINPUT34), .A2(KEYINPUT33), .ZN(n533) );
  NAND2_X1 U626 ( .A1(n534), .A2(n533), .ZN(n537) );
  NOR2_X1 U627 ( .A1(n535), .A2(n614), .ZN(n536) );
  NAND2_X1 U628 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U629 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n540) );
  NAND2_X1 U630 ( .A1(n576), .A2(KEYINPUT44), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n542), .B(KEYINPUT92), .ZN(n559) );
  INV_X1 U632 ( .A(n660), .ZN(n544) );
  NOR2_X1 U633 ( .A1(n544), .A2(n676), .ZN(n545) );
  XNOR2_X1 U634 ( .A(KEYINPUT104), .B(n545), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n551), .A2(n546), .ZN(n548) );
  XOR2_X1 U636 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n547) );
  NAND2_X1 U637 ( .A1(n571), .A2(n614), .ZN(n563) );
  INV_X1 U638 ( .A(n628), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n382), .A2(n427), .ZN(n549) );
  XNOR2_X2 U640 ( .A(n549), .B(KEYINPUT105), .ZN(n804) );
  INV_X1 U641 ( .A(n566), .ZN(n662) );
  AND2_X1 U642 ( .A1(n628), .A2(n426), .ZN(n667) );
  NAND2_X1 U643 ( .A1(n393), .A2(n667), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n550), .B(KEYINPUT31), .ZN(n767) );
  INV_X1 U645 ( .A(n656), .ZN(n552) );
  NOR2_X1 U646 ( .A1(n662), .A2(n552), .ZN(n553) );
  AND2_X1 U647 ( .A1(n555), .A2(n554), .ZN(n769) );
  INV_X1 U648 ( .A(n769), .ZN(n627) );
  OR2_X1 U649 ( .A1(n555), .A2(n554), .ZN(n616) );
  AND2_X1 U650 ( .A1(n627), .A2(n616), .ZN(n673) );
  NAND2_X1 U651 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U652 ( .A(n560), .B(KEYINPUT91), .ZN(n573) );
  XNOR2_X1 U653 ( .A(KEYINPUT32), .B(KEYINPUT65), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n561), .B(KEYINPUT81), .ZN(n565) );
  INV_X1 U655 ( .A(n659), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n657), .A2(n567), .ZN(n562) );
  NOR2_X1 U657 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U658 ( .A(n565), .B(n564), .Z(n801) );
  XNOR2_X1 U659 ( .A(n566), .B(KEYINPUT106), .ZN(n602) );
  NAND2_X1 U660 ( .A1(n380), .A2(n567), .ZN(n569) );
  INV_X1 U661 ( .A(n568), .ZN(n657) );
  NOR2_X1 U662 ( .A1(n569), .A2(n657), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n726) );
  NAND2_X1 U664 ( .A1(n801), .A2(n726), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n578), .A2(KEYINPUT44), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U667 ( .A(KEYINPUT90), .ZN(n574) );
  OR2_X1 U668 ( .A1(n728), .A2(KEYINPUT44), .ZN(n577) );
  OR2_X1 U669 ( .A1(n578), .A2(n577), .ZN(n579) );
  BUF_X1 U670 ( .A(n362), .Z(n582) );
  INV_X1 U671 ( .A(n582), .ZN(n583) );
  NAND2_X1 U672 ( .A1(n583), .A2(KEYINPUT84), .ZN(n640) );
  INV_X1 U673 ( .A(n678), .ZN(n599) );
  OR2_X1 U674 ( .A1(n584), .A2(G900), .ZN(n587) );
  INV_X1 U675 ( .A(n585), .ZN(n586) );
  AND2_X1 U676 ( .A1(n587), .A2(n586), .ZN(n600) );
  INV_X1 U677 ( .A(n600), .ZN(n588) );
  AND2_X1 U678 ( .A1(n656), .A2(n588), .ZN(n589) );
  AND2_X1 U679 ( .A1(n605), .A2(n589), .ZN(n607) );
  INV_X1 U680 ( .A(KEYINPUT76), .ZN(n592) );
  XNOR2_X1 U681 ( .A(n592), .B(KEYINPUT38), .ZN(n593) );
  AND2_X1 U682 ( .A1(n607), .A2(n675), .ZN(n594) );
  INV_X1 U683 ( .A(n616), .ZN(n596) );
  INV_X1 U684 ( .A(KEYINPUT40), .ZN(n597) );
  NOR2_X1 U685 ( .A1(n600), .A2(n659), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n660), .A2(n601), .ZN(n613) );
  OR2_X1 U687 ( .A1(n380), .A2(n613), .ZN(n603) );
  INV_X1 U688 ( .A(KEYINPUT110), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n606), .B(KEYINPUT46), .ZN(n624) );
  AND2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n611) );
  AND2_X1 U691 ( .A1(n591), .A2(n609), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U693 ( .A(n612), .B(KEYINPUT109), .ZN(n799) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT36), .ZN(n618) );
  OR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n762) );
  NOR2_X1 U697 ( .A1(n762), .A2(n673), .ZN(n622) );
  NOR2_X1 U698 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n366), .ZN(n626) );
  INV_X1 U701 ( .A(KEYINPUT48), .ZN(n625) );
  OR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT43), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n631), .A2(n403), .ZN(n633) );
  INV_X1 U705 ( .A(KEYINPUT108), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n800) );
  INV_X1 U707 ( .A(n800), .ZN(n634) );
  AND2_X1 U708 ( .A1(n725), .A2(n634), .ZN(n635) );
  NAND2_X2 U709 ( .A1(n636), .A2(n635), .ZN(n646) );
  XNOR2_X2 U710 ( .A(n646), .B(KEYINPUT87), .ZN(n701) );
  BUF_X2 U711 ( .A(n701), .Z(n710) );
  NOR2_X1 U712 ( .A1(n710), .A2(KEYINPUT85), .ZN(n638) );
  XNOR2_X1 U713 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n643) );
  INV_X1 U714 ( .A(n643), .ZN(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n645) );
  INV_X1 U717 ( .A(KEYINPUT85), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n641), .A2(KEYINPUT84), .ZN(n642) );
  OR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n655) );
  INV_X1 U721 ( .A(n646), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n647), .A2(KEYINPUT2), .ZN(n711) );
  INV_X1 U723 ( .A(n711), .ZN(n648) );
  INV_X1 U724 ( .A(KEYINPUT84), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n582), .A2(n649), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n710), .A2(KEYINPUT85), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n691) );
  XNOR2_X1 U730 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U734 ( .A(KEYINPUT49), .B(n661), .Z(n663) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U736 ( .A(KEYINPUT114), .B(n664), .Z(n665) );
  NOR2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n668) );
  OR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U739 ( .A(n670), .B(n669), .Z(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(KEYINPUT33), .ZN(n692) );
  INV_X1 U741 ( .A(n673), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U746 ( .A1(n692), .A2(n682), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n685), .B(KEYINPUT116), .ZN(n686) );
  XNOR2_X1 U749 ( .A(KEYINPUT52), .B(n686), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U751 ( .A(n689), .B(KEYINPUT117), .ZN(n690) );
  NAND2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U754 ( .A(KEYINPUT118), .B(n694), .Z(n695) );
  NOR2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U756 ( .A1(n795), .A2(n697), .ZN(n699) );
  XNOR2_X1 U757 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n698) );
  INV_X1 U758 ( .A(KEYINPUT2), .ZN(n700) );
  NAND2_X1 U759 ( .A1(n700), .A2(KEYINPUT86), .ZN(n702) );
  INV_X1 U760 ( .A(n701), .ZN(n794) );
  INV_X1 U761 ( .A(n702), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n794), .A2(n703), .ZN(n705) );
  NAND2_X1 U763 ( .A1(n708), .A2(KEYINPUT86), .ZN(n704) );
  NAND2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U765 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n714), .A2(n362), .ZN(n715) );
  INV_X1 U770 ( .A(KEYINPUT64), .ZN(n716) );
  NAND2_X1 U771 ( .A1(n750), .A2(G472), .ZN(n721) );
  XOR2_X1 U772 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n718) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X2 U774 ( .A1(n722), .A2(n754), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(G57) );
  XNOR2_X1 U776 ( .A(n725), .B(G134), .ZN(G36) );
  XNOR2_X1 U777 ( .A(n726), .B(G110), .ZN(G12) );
  XOR2_X1 U778 ( .A(n381), .B(G131), .Z(G33) );
  XOR2_X1 U779 ( .A(n728), .B(G122), .Z(G24) );
  NAND2_X1 U780 ( .A1(n744), .A2(G217), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n729), .B(KEYINPUT123), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n732), .A2(n754), .ZN(G66) );
  NAND2_X1 U784 ( .A1(n744), .A2(G478), .ZN(n735) );
  XOR2_X1 U785 ( .A(n733), .B(KEYINPUT122), .Z(n734) );
  XNOR2_X1 U786 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n736), .A2(n754), .ZN(G63) );
  NAND2_X1 U788 ( .A1(n750), .A2(G475), .ZN(n740) );
  XOR2_X1 U789 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n737) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X2 U791 ( .A1(n741), .A2(n754), .ZN(n743) );
  XNOR2_X1 U792 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G60) );
  NAND2_X1 U794 ( .A1(n744), .A2(G469), .ZN(n748) );
  XOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n749), .A2(n754), .ZN(G54) );
  BUF_X1 U799 ( .A(n751), .Z(n753) );
  XOR2_X1 U800 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n752) );
  XNOR2_X1 U801 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n755) );
  XOR2_X1 U802 ( .A(G104), .B(KEYINPUT113), .Z(n757) );
  NAND2_X1 U803 ( .A1(n758), .A2(n596), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n757), .B(n756), .ZN(G6) );
  XOR2_X1 U805 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n760) );
  NAND2_X1 U806 ( .A1(n758), .A2(n769), .ZN(n759) );
  XNOR2_X1 U807 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U808 ( .A(G107), .B(n761), .ZN(G9) );
  XOR2_X1 U809 ( .A(G128), .B(KEYINPUT29), .Z(n764) );
  INV_X1 U810 ( .A(n762), .ZN(n765) );
  NAND2_X1 U811 ( .A1(n765), .A2(n769), .ZN(n763) );
  XNOR2_X1 U812 ( .A(n764), .B(n763), .ZN(G30) );
  NAND2_X1 U813 ( .A1(n765), .A2(n596), .ZN(n766) );
  XNOR2_X1 U814 ( .A(n766), .B(G146), .ZN(G48) );
  NAND2_X1 U815 ( .A1(n596), .A2(n770), .ZN(n768) );
  XNOR2_X1 U816 ( .A(G113), .B(n768), .ZN(G15) );
  NAND2_X1 U817 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n771), .B(G116), .ZN(G18) );
  XOR2_X1 U819 ( .A(G125), .B(n772), .Z(n773) );
  XNOR2_X1 U820 ( .A(n773), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U821 ( .A1(n582), .A2(n795), .ZN(n778) );
  NAND2_X1 U822 ( .A1(G224), .A2(G953), .ZN(n774) );
  XNOR2_X1 U823 ( .A(n774), .B(KEYINPUT124), .ZN(n775) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n775), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G898), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n787) );
  BUF_X1 U827 ( .A(n779), .Z(n780) );
  XOR2_X1 U828 ( .A(KEYINPUT125), .B(n781), .Z(n782) );
  XNOR2_X1 U829 ( .A(n780), .B(n782), .ZN(n783) );
  XNOR2_X1 U830 ( .A(n783), .B(G101), .ZN(n785) );
  NOR2_X1 U831 ( .A1(n795), .A2(G898), .ZN(n784) );
  NOR2_X1 U832 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U833 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U834 ( .A(KEYINPUT126), .B(n788), .ZN(G69) );
  XNOR2_X1 U835 ( .A(n391), .B(n789), .ZN(n793) );
  XNOR2_X1 U836 ( .A(n793), .B(G227), .ZN(n791) );
  NAND2_X1 U837 ( .A1(G900), .A2(n791), .ZN(n792) );
  NAND2_X1 U838 ( .A1(n792), .A2(G953), .ZN(n798) );
  XNOR2_X1 U839 ( .A(n794), .B(n793), .ZN(n796) );
  NAND2_X1 U840 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U841 ( .A1(n798), .A2(n797), .ZN(G72) );
  XOR2_X1 U842 ( .A(G143), .B(n799), .Z(G45) );
  XOR2_X1 U843 ( .A(G140), .B(n800), .Z(G42) );
  XNOR2_X1 U844 ( .A(G119), .B(n801), .ZN(G21) );
  XNOR2_X1 U845 ( .A(G137), .B(KEYINPUT127), .ZN(n803) );
  XNOR2_X1 U846 ( .A(n803), .B(n802), .ZN(G39) );
  XOR2_X1 U847 ( .A(G101), .B(n804), .Z(n805) );
  XNOR2_X1 U848 ( .A(KEYINPUT112), .B(n805), .ZN(G3) );
endmodule

