//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n219), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G50), .B2(G226), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n218), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n216), .B1(new_n230), .B2(new_n211), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n214), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT67), .Z(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G226), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G232), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G41), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(G274), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n269), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G87), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n266), .A2(new_n278), .A3(KEYINPUT76), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT76), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n255), .B1(new_n274), .B2(new_n275), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n265), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n266), .A2(new_n278), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT16), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT7), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n272), .A2(new_n273), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n228), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G58), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n228), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n296), .B2(new_n201), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G159), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n288), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT7), .B1(new_n292), .B2(new_n208), .ZN(new_n302));
  NOR4_X1   g0102(.A1(new_n272), .A2(new_n273), .A3(new_n289), .A4(G20), .ZN(new_n303));
  OAI21_X1  g0103(.A(G68), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n300), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(KEYINPUT16), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n209), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n301), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G13), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n310), .A2(new_n208), .A3(G1), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT71), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n307), .B2(new_n209), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n208), .A2(G1), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n314), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n287), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT18), .B1(new_n287), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT77), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n309), .A2(new_n321), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n279), .A2(new_n328), .A3(new_n283), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n266), .A2(new_n278), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT17), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  AND4_X1   g0133(.A1(KEYINPUT17), .A2(new_n332), .A3(new_n309), .A4(new_n321), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n326), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  INV_X1    g0136(.A(new_n332), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n322), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n327), .A2(KEYINPUT17), .A3(new_n332), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT77), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n325), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n290), .A2(G222), .A3(new_n268), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT70), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n290), .A2(G1698), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n267), .B1(new_n219), .B2(new_n290), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n277), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n260), .A2(new_n262), .ZN(new_n348));
  INV_X1    g0148(.A(G41), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n264), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n255), .A2(new_n257), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G226), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n280), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n320), .A2(G50), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n311), .A2(new_n202), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n203), .A2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  INV_X1    g0159(.A(new_n298), .ZN(new_n360));
  INV_X1    g0160(.A(G33), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT72), .B1(new_n361), .B2(G20), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(new_n208), .A3(G33), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n358), .B1(new_n359), .B2(new_n360), .C1(new_n365), .C2(new_n313), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n318), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n357), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n347), .A2(new_n285), .A3(new_n351), .A4(new_n353), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n355), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT73), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n372), .A3(new_n368), .A4(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(new_n313), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT15), .B(G87), .Z(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n365), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n308), .A2(new_n319), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(new_n308), .B1(G77), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n311), .A2(new_n219), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n352), .A2(G244), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n290), .A2(G232), .A3(new_n268), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n385), .B1(new_n221), .B2(new_n290), .C1(new_n345), .C2(new_n229), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n350), .B(new_n384), .C1(new_n386), .C2(new_n277), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(G169), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n285), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n371), .A2(new_n373), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n347), .A2(G190), .A3(new_n351), .A4(new_n353), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT9), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n368), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n354), .A2(G200), .B1(new_n398), .B2(KEYINPUT10), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n368), .A2(new_n395), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n402), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n397), .A2(new_n399), .A3(new_n404), .A4(new_n400), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n387), .A2(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n383), .B(new_n406), .C1(new_n328), .C2(new_n387), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n393), .A2(new_n403), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n341), .B1(new_n408), .B2(KEYINPUT75), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT75), .B1(new_n410), .B2(new_n392), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n290), .B1(G232), .B2(new_n268), .ZN(new_n412));
  NOR2_X1   g0212(.A1(G226), .A2(G1698), .ZN(new_n413));
  INV_X1    g0213(.A(G97), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n412), .A2(new_n413), .B1(new_n361), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n350), .B1(new_n415), .B2(new_n277), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT13), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n352), .A2(G238), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n379), .A2(G68), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n312), .A2(KEYINPUT12), .A3(G68), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT12), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n311), .B2(new_n228), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n298), .A2(G50), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n427), .B1(new_n208), .B2(G68), .C1(new_n365), .C2(new_n219), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n318), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT11), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(KEYINPUT11), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n421), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n419), .A2(new_n420), .A3(new_n330), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n419), .A2(new_n420), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT14), .B1(new_n436), .B2(new_n280), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(G179), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n432), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n411), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n409), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n208), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT22), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT22), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n290), .A2(new_n448), .A3(new_n208), .A4(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n208), .A2(G107), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT23), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT24), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n450), .A2(KEYINPUT24), .A3(new_n451), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n308), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n319), .A2(G13), .B1(new_n256), .B2(G33), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n318), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n311), .A2(new_n221), .ZN(new_n463));
  XOR2_X1   g0263(.A(new_n463), .B(KEYINPUT25), .Z(new_n464));
  AND3_X1   g0264(.A1(new_n458), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n259), .A2(G1), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n255), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n222), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n290), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n290), .A2(G250), .A3(new_n268), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n479), .B2(new_n277), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G274), .A3(new_n466), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n480), .A2(new_n481), .A3(new_n330), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n330), .A3(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(new_n483), .ZN(new_n486));
  AOI211_X1 g0286(.A(new_n486), .B(new_n472), .C1(new_n479), .C2(new_n277), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n485), .B(KEYINPUT86), .C1(new_n487), .C2(G200), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n465), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n458), .A2(new_n462), .A3(new_n464), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n487), .A2(G169), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n285), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n308), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n302), .B2(new_n303), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  AND2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n298), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n495), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n318), .A2(new_n414), .A3(new_n460), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n311), .A2(new_n414), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT78), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G257), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n483), .B1(new_n471), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n277), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n277), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(KEYINPUT79), .A3(new_n277), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n508), .B(new_n519), .C1(new_n524), .C2(new_n328), .ZN(new_n525));
  INV_X1    g0325(.A(new_n510), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n517), .A2(KEYINPUT79), .A3(new_n277), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT79), .B1(new_n517), .B2(new_n277), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n285), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n518), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n280), .ZN(new_n531));
  INV_X1    g0331(.A(new_n505), .ZN(new_n532));
  INV_X1    g0332(.A(new_n507), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n496), .A2(new_n503), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n495), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n229), .A2(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n220), .A2(G1698), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n272), .C2(new_n273), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n277), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n264), .A2(new_n259), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n256), .A2(G45), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n255), .A2(G250), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n255), .B1(new_n539), .B2(new_n540), .ZN(new_n549));
  INV_X1    g0349(.A(new_n546), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n549), .A2(new_n543), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n312), .A2(new_n376), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n362), .A2(new_n364), .A3(G97), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n208), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n414), .A3(new_n221), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT80), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n290), .A2(new_n208), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n564), .A3(new_n560), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n556), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n553), .B1(new_n566), .B2(new_n308), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n308), .B(KEYINPUT71), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(KEYINPUT82), .A3(G87), .A4(new_n459), .ZN(new_n569));
  OAI211_X1 g0369(.A(G87), .B(new_n459), .C1(new_n315), .C2(new_n317), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n548), .A2(new_n552), .A3(new_n567), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(new_n308), .ZN(new_n575));
  INV_X1    g0375(.A(new_n553), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n376), .A3(new_n459), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n567), .A2(KEYINPUT81), .A3(new_n577), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n542), .A2(G179), .A3(new_n544), .A4(new_n546), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n551), .B2(new_n280), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n525), .A2(new_n536), .A3(new_n574), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n273), .ZN(new_n586));
  OR2_X1    g0386(.A1(KEYINPUT83), .A2(G303), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT3), .A2(G33), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT83), .A2(G303), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n277), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n277), .B1(new_n466), .B2(new_n482), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G270), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n483), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n311), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n459), .A2(G116), .A3(new_n495), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n307), .A2(new_n209), .B1(G20), .B2(new_n598), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n515), .B(new_n208), .C1(G33), .C2(new_n414), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(G169), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT84), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n597), .A2(new_n609), .A3(G169), .A4(new_n605), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n597), .A2(KEYINPUT21), .A3(G169), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n597), .A2(new_n285), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n605), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n597), .A2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(new_n605), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n615), .B(new_n616), .C1(new_n330), .C2(new_n597), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n494), .A2(new_n585), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n445), .A2(new_n619), .ZN(G372));
  NAND2_X1  g0420(.A1(new_n335), .A2(new_n340), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n441), .A2(new_n442), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n435), .A2(new_n391), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n325), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n403), .A2(new_n405), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n371), .A3(new_n373), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n536), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n518), .A2(G169), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n508), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(KEYINPUT87), .A3(new_n529), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n578), .A2(new_n583), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n574), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n567), .A2(KEYINPUT81), .A3(new_n577), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT81), .B1(new_n567), .B2(new_n577), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n549), .A2(new_n550), .A3(new_n285), .A4(new_n543), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(G169), .B2(new_n547), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n574), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n536), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n649));
  AOI22_X1  g0449(.A1(new_n633), .A2(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n489), .A2(new_n536), .A3(new_n525), .A4(new_n640), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n611), .A2(new_n614), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n639), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n445), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(new_n656), .ZN(G369));
  NOR2_X1   g0457(.A1(new_n310), .A2(G20), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .A3(G1), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT27), .B1(new_n659), .B2(G1), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n616), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n618), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n653), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n490), .A2(new_n664), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n489), .A2(new_n493), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT89), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n652), .A2(new_n664), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n489), .A2(KEYINPUT89), .A3(new_n493), .A4(new_n672), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n653), .A2(new_n665), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n675), .B2(new_n677), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n493), .A2(new_n664), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  INV_X1    g0485(.A(new_n212), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(G41), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n212), .A2(KEYINPUT90), .A3(new_n349), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n560), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n207), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n536), .A2(new_n634), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT87), .B1(new_n637), .B2(new_n529), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n640), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n648), .A2(new_n649), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n641), .B2(new_n633), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n639), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n525), .A2(new_n640), .A3(new_n536), .ZN(new_n703));
  INV_X1    g0503(.A(new_n488), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n458), .A2(new_n484), .A3(new_n462), .A4(new_n464), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n493), .A2(new_n614), .A3(new_n611), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n665), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n665), .B1(new_n655), .B2(new_n650), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT93), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT29), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n594), .A2(new_n483), .A3(new_n596), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n518), .A3(new_n480), .A4(new_n644), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT30), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n487), .A2(new_n719), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n285), .A3(new_n723), .A4(new_n547), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n665), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(KEYINPUT91), .A2(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT91), .B(KEYINPUT31), .Z(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n706), .A2(new_n652), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n536), .A2(new_n525), .A3(new_n574), .A4(new_n584), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n611), .A2(new_n614), .A3(new_n617), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .A4(new_n665), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n494), .A2(new_n618), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT92), .A3(new_n731), .A4(new_n665), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n729), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n718), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n693), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(new_n689), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n256), .B1(new_n658), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n209), .B1(G20), .B2(new_n280), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n208), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n328), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n208), .A2(new_n330), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n750), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n290), .B1(new_n751), .B2(new_n221), .C1(new_n559), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n285), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n749), .A2(new_n755), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n295), .B1(new_n757), .B2(new_n219), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n285), .A2(new_n328), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT95), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n759), .A2(new_n752), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(new_n759), .B2(new_n752), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n758), .B1(new_n764), .B2(G50), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n749), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G159), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n754), .B(new_n766), .C1(KEYINPUT32), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n767), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G97), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n759), .A2(new_n749), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(KEYINPUT32), .B2(new_n770), .C1(new_n228), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n757), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G311), .B1(new_n773), .B2(G294), .ZN(new_n779));
  INV_X1    g0579(.A(new_n753), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G303), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n779), .A2(new_n292), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G329), .B2(new_n769), .ZN(new_n783));
  INV_X1    g0583(.A(new_n751), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G283), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n764), .A2(G326), .ZN(new_n786));
  INV_X1    g0586(.A(new_n776), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  INV_X1    g0588(.A(new_n756), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(G322), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n748), .B1(new_n777), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n290), .A2(G355), .A3(new_n212), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n249), .A2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n686), .A2(new_n290), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n348), .A2(G50), .A3(new_n206), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n793), .B1(G116), .B2(new_n212), .C1(new_n794), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n747), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n669), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n746), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n746), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n669), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n671), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT97), .Z(G396));
  NOR2_X1   g0611(.A1(new_n391), .A2(new_n664), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n382), .A2(new_n664), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n407), .A2(new_n813), .B1(new_n389), .B2(new_n390), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n712), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n665), .B(new_n815), .C1(new_n655), .C2(new_n650), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n740), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n807), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n807), .B1(new_n816), .B2(new_n799), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n774), .B1(new_n221), .B2(new_n753), .C1(new_n823), .C2(new_n776), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G303), .B2(new_n764), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n751), .A2(new_n559), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n292), .B1(new_n757), .B2(new_n598), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G294), .C2(new_n789), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(new_n829), .C2(new_n768), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G150), .A2(new_n787), .B1(new_n789), .B2(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n757), .C1(new_n763), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT34), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n784), .A2(G68), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n202), .B2(new_n753), .C1(new_n837), .C2(new_n768), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n835), .A2(new_n292), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n773), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n295), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n830), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n747), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n747), .A2(new_n799), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n822), .B(new_n843), .C1(G77), .C2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n821), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NAND2_X1  g0648(.A1(new_n735), .A2(new_n737), .ZN(new_n849));
  OR2_X1    g0649(.A1(KEYINPUT102), .A2(KEYINPUT31), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n725), .B(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n816), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n327), .A2(new_n332), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n287), .A2(new_n322), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(new_n662), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n322), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n301), .A2(new_n306), .A3(new_n318), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n321), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n857), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n287), .A2(new_n861), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n854), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n859), .B1(new_n864), .B2(new_n856), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n341), .B2(new_n862), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n865), .B(KEYINPUT38), .C1(new_n341), .C2(new_n862), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(KEYINPUT98), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n341), .A2(new_n862), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT98), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT38), .A4(new_n865), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n432), .A2(new_n665), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n623), .A2(new_n664), .B1(new_n443), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n853), .A2(new_n870), .A3(new_n873), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n851), .B1(new_n735), .B2(new_n737), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n880), .A2(new_n816), .A3(new_n876), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT100), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(new_n859), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n338), .A2(new_n339), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n322), .B(new_n857), .C1(new_n325), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n859), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n882), .B1(new_n891), .B2(new_n869), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n878), .A2(new_n879), .B1(new_n881), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT92), .B1(new_n619), .B2(new_n665), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n732), .A2(new_n489), .A3(new_n493), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n895), .A2(new_n734), .A3(new_n585), .A4(new_n664), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n852), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n445), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n870), .A2(new_n873), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n815), .A3(new_n877), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n879), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n881), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(G330), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n445), .A2(G330), .A3(new_n897), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n898), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n631), .B1(new_n718), .B2(new_n445), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n622), .A2(new_n664), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n870), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n891), .A2(new_n913), .A3(new_n869), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n911), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n325), .A2(new_n662), .ZN(new_n916));
  INV_X1    g0716(.A(new_n812), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n876), .B1(new_n818), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n899), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n909), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n256), .B2(new_n658), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n598), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n209), .A2(new_n208), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(KEYINPUT35), .C2(new_n502), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  OAI21_X1  g0728(.A(G77), .B1(new_n295), .B2(new_n228), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n207), .A2(new_n929), .B1(G50), .B2(new_n228), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n310), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(G367));
  INV_X1    g0732(.A(new_n681), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n535), .A2(new_n664), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n525), .A2(new_n536), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n936));
  INV_X1    g0736(.A(new_n536), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n664), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT103), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n525), .A2(new_n939), .A3(new_n536), .A4(new_n934), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT42), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n681), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n936), .A2(new_n940), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n937), .B1(new_n946), .B2(new_n652), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n943), .B(new_n945), .C1(new_n947), .C2(new_n664), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n665), .B1(new_n567), .B2(new_n573), .ZN(new_n949));
  MUX2_X1   g0749(.A(new_n640), .B(new_n702), .S(new_n949), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT104), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT104), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n955), .A3(new_n951), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n953), .B2(new_n956), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(new_n679), .B2(new_n942), .ZN(new_n960));
  INV_X1    g0760(.A(new_n959), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n679), .A2(new_n942), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n689), .B(KEYINPUT41), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n679), .ZN(new_n966));
  INV_X1    g0766(.A(new_n683), .ZN(new_n967));
  NAND2_X1  g0767(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n968));
  OR2_X1    g0768(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n967), .A2(new_n942), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n683), .C2(new_n941), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT45), .B1(new_n683), .B2(new_n941), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n681), .A2(new_n942), .A3(new_n974), .A4(new_n682), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n966), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n680), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n671), .B1(new_n979), .B2(new_n681), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n933), .A2(new_n670), .A3(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n729), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n894), .B2(new_n896), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(G330), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n714), .A2(new_n982), .A3(new_n985), .A4(new_n717), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT106), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n973), .A2(new_n975), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n988), .A2(new_n679), .A3(new_n971), .A4(new_n970), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n710), .A2(new_n665), .B1(new_n712), .B2(KEYINPUT93), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n716), .B1(new_n990), .B2(KEYINPUT29), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(new_n985), .A4(new_n982), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n977), .A2(new_n987), .A3(new_n989), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n965), .B1(new_n994), .B2(new_n741), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n960), .B(new_n963), .C1(new_n995), .C2(new_n745), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n290), .B1(new_n751), .B2(new_n219), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G58), .A2(new_n780), .B1(new_n789), .B2(G150), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n840), .A2(new_n228), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n764), .B2(G143), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n202), .B2(new_n757), .C1(new_n833), .C2(new_n768), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(G159), .C2(new_n787), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n784), .A2(G97), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n292), .C1(new_n1007), .C2(new_n768), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n587), .A2(new_n589), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1009), .A2(new_n789), .B1(new_n778), .B2(G283), .ZN(new_n1010));
  INV_X1    g0810(.A(G294), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n776), .C1(new_n763), .C2(new_n829), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1008), .B(new_n1012), .C1(G107), .C2(new_n773), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT107), .B1(new_n753), .B2(new_n598), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT46), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n1005), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n747), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n950), .A2(new_n804), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n795), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n802), .B1(new_n212), .B2(new_n377), .C1(new_n238), .C2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n746), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n996), .A2(new_n1022), .ZN(G387));
  AND2_X1   g0823(.A1(new_n986), .A2(new_n743), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT113), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT113), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n741), .C2(new_n982), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n764), .A2(G322), .B1(G311), .B2(new_n787), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT111), .Z(new_n1029));
  AOI22_X1  g0829(.A1(G317), .A2(new_n789), .B1(new_n778), .B2(new_n1009), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT48), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n823), .B2(new_n840), .C1(new_n1011), .C2(new_n753), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n769), .A2(G326), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n292), .B1(new_n751), .B2(new_n598), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1006), .B1(new_n202), .B2(new_n756), .C1(new_n313), .C2(new_n776), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n840), .A2(new_n377), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n292), .B(new_n1040), .C1(new_n764), .C2(G159), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n228), .B2(new_n757), .C1(new_n219), .C2(new_n753), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(G150), .C2(new_n769), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT110), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n747), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n690), .B(new_n259), .C1(new_n228), .C2(new_n219), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT109), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n374), .A2(new_n202), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n795), .B1(new_n1047), .B2(new_n1049), .C1(new_n244), .C2(new_n348), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n290), .A2(new_n212), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(G107), .B2(new_n212), .C1(new_n690), .C2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n807), .B1(new_n1052), .B2(new_n802), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1045), .B(new_n1053), .C1(new_n678), .C2(new_n804), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n982), .A2(new_n745), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1027), .A2(new_n1056), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n977), .A2(new_n989), .A3(new_n745), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n942), .A2(new_n801), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n763), .A2(new_n1007), .B1(new_n829), .B2(new_n756), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n787), .A2(new_n1009), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n778), .A2(G294), .B1(new_n773), .B2(G116), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n753), .A2(new_n823), .B1(new_n751), .B2(new_n221), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n290), .B(new_n1064), .C1(G322), .C2(new_n769), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n763), .A2(new_n359), .B1(new_n832), .B2(new_n756), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT51), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n787), .B1(new_n778), .B2(new_n374), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1072), .A2(new_n292), .A3(new_n826), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n769), .A2(G143), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n753), .A2(new_n228), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n840), .A2(new_n219), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1066), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n747), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n802), .B1(new_n414), .B2(new_n212), .C1(new_n252), .C2(new_n1020), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1059), .A2(new_n746), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n977), .A2(new_n989), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n689), .B1(new_n1084), .B2(new_n986), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(KEYINPUT115), .A3(new_n994), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT115), .B1(new_n1085), .B2(new_n994), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1058), .B(new_n1083), .C1(new_n1087), .C2(new_n1088), .ZN(G390));
  INV_X1    g0889(.A(new_n445), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n632), .B(new_n905), .C1(new_n991), .C2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n984), .A2(G330), .A3(new_n815), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n876), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n853), .A2(G330), .A3(new_n877), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n641), .A2(new_n633), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n648), .A2(new_n649), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n664), .B1(new_n709), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n812), .B1(new_n1099), .B2(new_n815), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n740), .A2(new_n815), .A3(new_n877), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n664), .B1(new_n701), .B2(new_n709), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n814), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n812), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n880), .A2(new_n739), .A3(new_n816), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1106), .C1(new_n1107), .C2(new_n877), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1091), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n911), .C1(new_n1100), .C2(new_n876), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT116), .B1(new_n918), .B2(new_n910), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n912), .A4(new_n914), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n891), .A2(new_n869), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n911), .B(new_n1114), .C1(new_n1106), .C2(new_n876), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1094), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1103), .A3(new_n1115), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1109), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n877), .B1(new_n853), .B2(G330), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n738), .A2(new_n739), .A3(new_n816), .A4(new_n876), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n917), .B1(new_n711), .B2(new_n814), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1100), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n908), .B(new_n905), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1113), .A2(new_n1103), .A3(new_n1115), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1094), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1120), .A2(new_n1129), .A3(new_n743), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1120), .A2(new_n1129), .A3(KEYINPUT117), .A4(new_n743), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n912), .A2(new_n799), .A3(new_n914), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n845), .A2(new_n374), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n290), .B1(new_n764), .B2(G283), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n414), .B2(new_n757), .C1(new_n221), .C2(new_n776), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n753), .A2(new_n559), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n836), .B1(new_n598), .B2(new_n756), .C1(new_n1011), .C2(new_n768), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1077), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n751), .A2(new_n202), .B1(new_n768), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n764), .A2(G128), .B1(G132), .B2(new_n789), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT54), .B(G143), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n778), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n787), .A2(G137), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1145), .A2(new_n290), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1144), .B(new_n1149), .C1(G159), .C2(new_n773), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n753), .A2(new_n359), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1142), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n807), .B(new_n1137), .C1(new_n1154), .C2(new_n747), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1135), .A2(new_n745), .B1(new_n1136), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1134), .A2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n403), .A2(new_n370), .A3(new_n405), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT121), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT121), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n403), .A2(new_n1161), .A3(new_n370), .A4(new_n405), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n368), .A2(new_n857), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1169), .A3(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n903), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n893), .A2(G330), .A3(new_n1173), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1175), .A2(new_n921), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n921), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1091), .B1(new_n1135), .B2(new_n1109), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1158), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1173), .B1(new_n893), .B2(G330), .ZN(new_n1182));
  AND4_X1   g0982(.A1(G330), .A2(new_n901), .A3(new_n902), .A4(new_n1173), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n922), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1175), .A2(new_n1176), .A3(new_n921), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1091), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1120), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1178), .A2(KEYINPUT122), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1189), .A3(KEYINPUT57), .A4(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1181), .A2(new_n1191), .A3(new_n743), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1174), .A2(new_n799), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n776), .A2(new_n837), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1146), .ZN(new_n1195));
  INV_X1    g0995(.A(G128), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1195), .A2(new_n753), .B1(new_n1196), .B2(new_n756), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n1143), .B2(new_n763), .C1(new_n359), .C2(new_n840), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1194), .B(new_n1199), .C1(G137), .C2(new_n778), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G41), .B1(new_n769), .B2(G124), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G33), .B1(new_n784), .B2(G159), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n202), .B1(new_n272), .B2(G41), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n349), .B1(new_n753), .B2(new_n219), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1207), .B(new_n1002), .C1(G97), .C2(new_n787), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n292), .B1(new_n768), .B2(new_n823), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n756), .A2(new_n221), .B1(new_n751), .B2(new_n295), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n376), .C2(new_n778), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(new_n598), .C2(new_n763), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT58), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1205), .A2(new_n1206), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n747), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n844), .A2(new_n202), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1193), .A2(new_n746), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1219), .B2(new_n745), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1192), .A2(new_n1220), .ZN(G375));
  OAI21_X1  g1021(.A(new_n746), .B1(G68), .B2(new_n845), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n753), .A2(new_n414), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n290), .B1(new_n764), .B2(G294), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n221), .B2(new_n757), .C1(new_n598), .C2(new_n776), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G303), .C2(new_n769), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1040), .B1(G77), .B2(new_n784), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n823), .C2(new_n756), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT123), .Z(new_n1229));
  AOI22_X1  g1029(.A1(new_n784), .A2(G58), .B1(new_n773), .B2(G50), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n1196), .B2(new_n768), .C1(new_n776), .C2(new_n1195), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G137), .B2(new_n789), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n290), .B1(new_n763), .B2(new_n837), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G150), .B2(new_n778), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(new_n832), .C2(new_n753), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n748), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1222), .B(new_n1236), .C1(new_n799), .C2(new_n876), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n745), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n964), .B1(new_n1238), .B2(new_n1188), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1240), .B2(new_n1109), .ZN(G381));
  INV_X1    g1041(.A(new_n1083), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1085), .A2(new_n994), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT115), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1245), .B2(new_n1086), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(new_n996), .A3(new_n1022), .A4(new_n1058), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G381), .A2(G384), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1247), .A2(G396), .A3(G393), .A4(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1130), .A2(new_n1156), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1220), .A3(new_n1192), .A4(new_n1250), .ZN(G407));
  NOR2_X1   g1051(.A1(new_n1249), .A2(new_n663), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1192), .A2(new_n1220), .A3(new_n1250), .ZN(new_n1253));
  OAI21_X1  g1053(.A(G213), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G378), .A2(new_n1192), .A3(new_n1220), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1187), .A2(new_n745), .A3(new_n1190), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1189), .A2(new_n1219), .A3(new_n964), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1217), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1250), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1238), .B2(new_n1188), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1102), .A2(new_n1091), .A3(new_n1108), .A4(KEYINPUT60), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n743), .A3(new_n1126), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1239), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n847), .A2(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n847), .A2(KEYINPUT125), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1257), .A2(G2897), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n847), .A4(new_n1239), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1263), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  INV_X1    g1079(.A(G396), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G390), .A2(G387), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1247), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1247), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1278), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1257), .B(new_n1288), .C1(new_n1258), .C2(new_n1262), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT63), .B1(new_n1289), .B2(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1288), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1263), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT126), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1287), .A2(new_n1290), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1263), .A2(new_n1297), .A3(new_n1291), .ZN(new_n1298));
  XOR2_X1   g1098(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1263), .B2(new_n1276), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1263), .B2(new_n1291), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1247), .A2(new_n1283), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1247), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1296), .B1(new_n1302), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1250), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1258), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1307), .B(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1288), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1307), .B1(new_n1258), .B2(new_n1309), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1306), .B2(new_n1305), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1291), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(G402));
endmodule


