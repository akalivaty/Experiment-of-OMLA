//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AND2_X1   g0007(.A1(G87), .A2(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n208), .B(new_n213), .C1(G116), .C2(G270), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n203), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n207), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n222), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT64), .ZN(G361));
  XOR2_X1   g0031(.A(G226), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G222), .B2(G1698), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G77), .B2(new_n254), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n257), .B(G274), .C1(G41), .C2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n250), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G169), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n204), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  INV_X1    g0069(.A(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n265), .B1(new_n266), .B2(new_n268), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n226), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n257), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n201), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n264), .B(new_n281), .C1(G179), .C2(new_n262), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT10), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(G200), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(KEYINPUT70), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT9), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n281), .A2(new_n288), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n281), .A2(new_n288), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n289), .A3(KEYINPUT9), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n284), .B1(new_n296), .B2(new_n262), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n286), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n285), .B(new_n297), .C1(new_n292), .C2(new_n294), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n282), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  INV_X1    g0102(.A(new_n258), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n259), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n304), .A2(new_n211), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n250), .A2(G238), .A3(new_n260), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n302), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n250), .B1(new_n312), .B2(new_n314), .ZN(new_n321));
  NOR4_X1   g0121(.A1(new_n321), .A2(KEYINPUT13), .A3(new_n318), .A4(new_n303), .ZN(new_n322));
  OAI21_X1  g0122(.A(G200), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n307), .A2(new_n311), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n313), .B1(new_n324), .B2(new_n254), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n258), .B(new_n319), .C1(new_n325), .C2(new_n250), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n317), .A2(new_n302), .A3(new_n319), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G190), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n276), .A2(G68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT12), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n279), .B2(new_n203), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n209), .B2(new_n271), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n274), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT11), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(KEYINPUT11), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n323), .A2(new_n329), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT71), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n323), .A2(new_n329), .A3(KEYINPUT71), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n320), .B2(new_n322), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n327), .A2(new_n328), .A3(G179), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(G169), .C1(new_n320), .C2(new_n322), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n340), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n301), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G20), .A2(G77), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n356), .B1(new_n358), .B2(new_n271), .C1(new_n268), .C2(new_n269), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n274), .B1(G77), .B2(new_n276), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n278), .A2(G77), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G238), .A2(G1698), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n254), .B(new_n364), .C1(new_n310), .C2(G1698), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n316), .C1(G107), .C2(new_n254), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n258), .B1(new_n261), .B2(new_n210), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT67), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT67), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n258), .C1(new_n261), .C2(new_n210), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n263), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n363), .B(new_n372), .C1(G179), .C2(new_n371), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n254), .B2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n254), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n305), .A2(new_n309), .ZN(new_n379));
  INV_X1    g0179(.A(new_n377), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(KEYINPUT72), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G68), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n202), .A2(new_n203), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n267), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n304), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n309), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT73), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n380), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n203), .B1(new_n395), .B2(new_n375), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n391), .B1(new_n396), .B2(new_n388), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n274), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n269), .A2(new_n278), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n276), .B2(new_n269), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n251), .A2(new_n306), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n259), .A2(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n305), .A2(new_n401), .A3(new_n309), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n316), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n250), .A2(new_n260), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n303), .B1(new_n407), .B2(G232), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(new_n296), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n250), .B1(new_n403), .B2(new_n404), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n258), .B1(new_n261), .B2(new_n310), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(KEYINPUT74), .A3(new_n413), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n398), .A2(new_n400), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n417), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT74), .B1(new_n409), .B2(new_n413), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n398), .A4(new_n400), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n398), .A2(new_n400), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n263), .B1(new_n406), .B2(new_n408), .ZN(new_n426));
  INV_X1    g0226(.A(G179), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n411), .A2(new_n412), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT18), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n432), .B(new_n429), .C1(new_n398), .C2(new_n400), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n420), .B(new_n424), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n371), .A2(new_n296), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n371), .A2(G200), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n360), .A3(new_n362), .A4(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n355), .A2(new_n373), .A3(new_n435), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n210), .A2(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n305), .A3(new_n309), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n305), .A2(new_n309), .A3(G250), .A4(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n441), .A2(new_n305), .A3(new_n309), .A4(KEYINPUT4), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n316), .ZN(new_n449));
  XOR2_X1   g0249(.A(KEYINPUT5), .B(G41), .Z(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G274), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n452), .B1(new_n227), .B2(new_n249), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(G257), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT75), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n449), .A2(new_n460), .A3(new_n457), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(G200), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n449), .A2(G190), .A3(new_n457), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n464), .A2(new_n211), .A3(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(G97), .B(G107), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(new_n270), .B1(new_n209), .B2(new_n268), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n395), .B2(new_n375), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n274), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n278), .A2(G97), .ZN(new_n472));
  INV_X1    g0272(.A(new_n274), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n257), .A2(G33), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n473), .A2(new_n278), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(G97), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n463), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n254), .A2(new_n270), .A3(G68), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT19), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n271), .B2(new_n211), .ZN(new_n481));
  NOR3_X1   g0281(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n313), .B2(KEYINPUT19), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n274), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n475), .A2(new_n357), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n358), .A2(new_n279), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n257), .A2(G45), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n250), .A2(G250), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n453), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n219), .A2(new_n306), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n210), .A2(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n254), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n491), .B1(new_n496), .B2(new_n316), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n427), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n250), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n263), .B1(new_n499), .B2(new_n491), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(G190), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n484), .A2(new_n274), .B1(new_n358), .B2(new_n279), .ZN(new_n503));
  OAI21_X1  g0303(.A(G200), .B1(new_n499), .B2(new_n491), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n475), .A2(G87), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n449), .A2(G179), .A3(new_n457), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(new_n250), .C1(new_n450), .C2(new_n489), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n455), .A2(G274), .A3(new_n452), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n316), .B2(new_n448), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n508), .B1(new_n512), .B2(new_n263), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n471), .A2(new_n476), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(G250), .A2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n212), .A2(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n305), .A2(new_n516), .A3(new_n309), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G294), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n316), .A2(new_n520), .B1(new_n456), .B2(G264), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n296), .A3(new_n510), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n316), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n456), .A2(G264), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n523), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n525), .B2(G200), .ZN(new_n526));
  AND4_X1   g0326(.A1(new_n270), .A2(new_n305), .A3(new_n309), .A4(G87), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT78), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT77), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(KEYINPUT22), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(KEYINPUT77), .A3(KEYINPUT78), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n527), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n270), .B2(G107), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT23), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n270), .A2(G33), .A3(G116), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n537), .B(KEYINPUT23), .C1(new_n270), .C2(G107), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n533), .A2(new_n534), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n305), .A2(new_n309), .A3(new_n270), .A4(G87), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n529), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n536), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n536), .A2(new_n543), .A3(KEYINPUT24), .A4(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n274), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n475), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n278), .A2(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT25), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n526), .A2(new_n551), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n478), .A2(new_n507), .A3(new_n515), .A4(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT80), .B1(new_n525), .B2(new_n263), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n521), .A2(new_n510), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT80), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(G169), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n525), .A2(G179), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n454), .B1(G270), .B2(new_n456), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n316), .B1(new_n254), .B2(G303), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n306), .A2(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G264), .A2(G1698), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n305), .A2(new_n309), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n566), .A2(new_n569), .A3(KEYINPUT76), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT76), .ZN(new_n571));
  INV_X1    g0371(.A(G303), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n250), .B1(new_n379), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n254), .A2(new_n567), .A3(new_n568), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n565), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n473), .A2(G116), .A3(new_n278), .A4(new_n474), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n273), .A2(new_n226), .B1(G20), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n445), .B(new_n270), .C1(G33), .C2(new_n211), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI221_X1 g0382(.A(new_n577), .B1(G116), .B2(new_n278), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(G169), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n576), .A2(G200), .ZN(new_n587));
  INV_X1    g0387(.A(new_n583), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT76), .B1(new_n566), .B2(new_n569), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(new_n571), .A3(new_n574), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G190), .A3(new_n565), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n576), .A2(KEYINPUT21), .A3(new_n583), .A4(G169), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n583), .A2(G179), .A3(new_n591), .A4(new_n565), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n586), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n556), .A2(new_n564), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n440), .A2(new_n597), .ZN(G372));
  NOR2_X1   g0398(.A1(new_n431), .A2(new_n433), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n345), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n353), .B1(new_n601), .B2(new_n373), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n420), .A2(new_n424), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n290), .A2(new_n291), .A3(new_n287), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT9), .B1(new_n293), .B2(new_n289), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n298), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n285), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n295), .A2(new_n286), .A3(new_n298), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n282), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n556), .A2(KEYINPUT81), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n586), .A2(new_n594), .A3(new_n595), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n562), .A2(new_n563), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n586), .A2(KEYINPUT82), .A3(new_n594), .A4(new_n595), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n462), .A2(new_n477), .B1(new_n513), .B2(new_n514), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT81), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n507), .A4(new_n555), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n501), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n513), .A2(new_n514), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n507), .A3(KEYINPUT26), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n513), .A2(new_n501), .A3(new_n506), .A4(new_n514), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n626), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n440), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n614), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(G13), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n257), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n588), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n596), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n618), .A2(new_n620), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n645), .ZN(new_n648));
  INV_X1    g0448(.A(G330), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n619), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n563), .A2(new_n643), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n555), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n619), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n651), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n586), .A2(new_n594), .A3(new_n595), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n643), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n223), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G1), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n482), .A2(new_n578), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n229), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n633), .A2(new_n644), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT86), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT29), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n643), .B1(new_n625), .B2(new_n632), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT86), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n629), .A2(new_n676), .A3(new_n630), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT87), .B1(new_n629), .B2(new_n630), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n627), .A2(new_n507), .A3(new_n679), .A4(KEYINPUT26), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n675), .A2(new_n677), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n657), .A2(new_n619), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n506), .A3(new_n622), .A4(new_n555), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n683), .A3(new_n501), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n671), .B1(new_n684), .B2(new_n644), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n674), .A2(new_n686), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n507), .A2(new_n478), .A3(new_n515), .A4(new_n555), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n564), .A2(new_n596), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n644), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n591), .A2(new_n497), .A3(new_n521), .A4(new_n565), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT84), .B1(new_n691), .B2(new_n508), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT30), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT84), .B(new_n694), .C1(new_n691), .C2(new_n508), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n512), .A2(new_n525), .ZN(new_n696));
  INV_X1    g0496(.A(new_n497), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n427), .A3(new_n697), .A4(new_n576), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n643), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n690), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT85), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n707), .A3(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n687), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n667), .B1(new_n710), .B2(G1), .ZN(G364));
  AOI21_X1  g0511(.A(new_n664), .B1(G45), .B2(new_n637), .ZN(new_n712));
  INV_X1    g0512(.A(new_n650), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n648), .A2(new_n649), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n712), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n226), .B1(G20), .B2(new_n263), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n270), .A2(new_n296), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n427), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n270), .A2(G190), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G179), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(G322), .A2(new_n724), .B1(new_n728), .B2(G329), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n427), .A2(new_n410), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n725), .ZN(new_n731));
  XOR2_X1   g0531(.A(KEYINPUT33), .B(G317), .Z(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n410), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n379), .B1(new_n735), .B2(new_n572), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n721), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(G326), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n725), .A2(new_n722), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n726), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n733), .B(new_n742), .C1(G294), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G283), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n725), .A2(new_n734), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n731), .ZN(new_n749));
  INV_X1    g0549(.A(new_n735), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G68), .A2(new_n749), .B1(new_n750), .B2(G87), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n202), .B2(new_n723), .ZN(new_n752));
  INV_X1    g0552(.A(G159), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n727), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT92), .B(KEYINPUT32), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n744), .A2(G97), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n747), .A2(new_n469), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n379), .B(new_n759), .C1(G50), .C2(new_n738), .ZN(new_n760));
  INV_X1    g0560(.A(new_n754), .ZN(new_n761));
  INV_X1    g0561(.A(new_n741), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(new_n755), .B1(G77), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n757), .A2(new_n758), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n748), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n648), .A2(new_n719), .B1(new_n720), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(G355), .B(KEYINPUT89), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n223), .A3(new_n254), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G116), .B2(new_n223), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT90), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n661), .A2(new_n254), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n247), .B2(G45), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G45), .B2(new_n229), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT91), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n719), .A2(new_n720), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n716), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n715), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT93), .ZN(G396));
  OR2_X1    g0581(.A1(new_n373), .A2(new_n643), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n363), .A2(new_n643), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n438), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n373), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n717), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n758), .B1(new_n578), .B2(new_n741), .C1(new_n572), .C2(new_n737), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G283), .B2(new_n749), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n254), .B1(new_n750), .B2(G107), .ZN(new_n790));
  INV_X1    g0590(.A(new_n747), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G294), .A2(new_n724), .B1(new_n791), .B2(G87), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n728), .A2(G311), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n789), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n724), .B1(new_n762), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n737), .C1(new_n266), .C2(new_n731), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n254), .B1(new_n735), .B2(new_n201), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n747), .A2(new_n203), .B1(new_n727), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(G58), .C2(new_n744), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  OAI21_X1  g0603(.A(new_n794), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n720), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n720), .A2(new_n717), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n209), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n787), .A2(new_n712), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT86), .B1(new_n633), .B2(new_n644), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n669), .B(new_n643), .C1(new_n625), .C2(new_n632), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n786), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT95), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n672), .A2(new_n813), .A3(new_n812), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n672), .B2(new_n812), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(new_n709), .Z(new_n817));
  OAI21_X1  g0617(.A(new_n808), .B1(new_n817), .B2(new_n712), .ZN(G384));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n687), .A2(new_n819), .A3(new_n440), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n687), .B2(new_n440), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n614), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT96), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n373), .A2(new_n643), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n633), .A2(new_n644), .A3(new_n812), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT95), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n672), .A2(new_n813), .A3(new_n812), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n352), .A2(new_n643), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n345), .A2(new_n353), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n345), .B2(new_n353), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n824), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n782), .B1(new_n814), .B2(new_n815), .ZN(new_n836));
  INV_X1    g0636(.A(new_n834), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(KEYINPUT96), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n388), .B1(new_n382), .B2(G68), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n473), .B1(new_n839), .B2(KEYINPUT16), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT16), .B2(new_n839), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n641), .B1(new_n841), .B2(new_n400), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n599), .B2(new_n604), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n841), .A2(new_n400), .B1(new_n429), .B2(new_n641), .ZN(new_n844));
  INV_X1    g0644(.A(new_n418), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n641), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n425), .B1(new_n430), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n418), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n835), .A2(new_n838), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n599), .A2(new_n641), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT97), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n425), .A2(new_n847), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n398), .A2(new_n400), .B1(new_n429), .B2(new_n641), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n845), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n434), .A2(new_n862), .B1(new_n850), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n860), .B1(new_n865), .B2(KEYINPUT38), .ZN(new_n866));
  MUX2_X1   g0666(.A(new_n860), .B(new_n866), .S(new_n854), .Z(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n867), .B2(new_n858), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n353), .A2(new_n643), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n856), .A2(new_n857), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n823), .B(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n843), .A2(KEYINPUT97), .A3(new_n851), .A4(KEYINPUT38), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT40), .B(new_n873), .C1(new_n866), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n830), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n354), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n786), .B1(new_n877), .B2(new_n831), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT100), .B1(new_n700), .B2(new_n701), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT100), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n880), .B(KEYINPUT31), .C1(new_n699), .C2(new_n643), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n690), .A2(new_n703), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n874), .A2(new_n852), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(new_n884), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n703), .B(new_n690), .C1(new_n879), .C2(new_n881), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n878), .C1(new_n874), .C2(new_n852), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n885), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n866), .A2(new_n874), .ZN(new_n898));
  INV_X1    g0698(.A(new_n884), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT40), .A4(new_n873), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT101), .B1(new_n893), .B2(new_n887), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n900), .B(G330), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n440), .A2(G330), .A3(new_n892), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n897), .A2(new_n440), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n872), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n257), .B2(new_n637), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT35), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n228), .B1(new_n467), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(G116), .C1(new_n908), .C2(new_n467), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  OAI21_X1  g0711(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n912), .A2(new_n229), .B1(G50), .B2(new_n203), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(G1), .A3(new_n636), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n911), .A3(new_n914), .ZN(G367));
  NAND2_X1  g0715(.A1(new_n503), .A2(new_n505), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n643), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n507), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(new_n501), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n627), .A2(new_n643), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n514), .A2(new_n643), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n622), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n654), .A3(new_n658), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT42), .A3(new_n930), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n925), .A2(new_n927), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n515), .B1(new_n936), .B2(new_n619), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n644), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n921), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n655), .A2(new_n936), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n921), .A3(new_n940), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n939), .A2(new_n921), .A3(new_n940), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n946), .A2(new_n941), .B1(new_n655), .B2(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n662), .B(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n659), .A2(new_n656), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n950), .A2(new_n936), .A3(KEYINPUT44), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT44), .B1(new_n950), .B2(new_n936), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n950), .B2(new_n936), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n928), .A2(new_n659), .A3(new_n656), .A4(new_n955), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n655), .A2(KEYINPUT105), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n654), .B(new_n658), .Z(new_n964));
  NOR2_X1   g0764(.A1(new_n650), .A2(KEYINPUT106), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n710), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n961), .A2(new_n962), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n710), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n949), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n257), .B1(new_n637), .B2(G45), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n948), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n731), .A2(new_n753), .B1(new_n741), .B2(new_n201), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT107), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(new_n254), .C1(new_n202), .C2(new_n735), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n727), .A2(new_n796), .ZN(new_n978));
  INV_X1    g0778(.A(new_n744), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n203), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G143), .A2(new_n738), .B1(new_n724), .B2(G150), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n209), .B2(new_n747), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT108), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n723), .A2(new_n572), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n254), .B1(new_n762), .B2(G283), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n740), .B2(new_n737), .C1(new_n987), .C2(new_n727), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n985), .B(new_n988), .C1(G107), .C2(new_n744), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n791), .A2(G97), .ZN(new_n990));
  INV_X1    g0790(.A(G294), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(new_n731), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n735), .A2(new_n578), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n984), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n720), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n918), .A2(new_n719), .A3(new_n919), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n777), .B1(new_n223), .B2(new_n358), .C1(new_n239), .C2(new_n772), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n997), .A2(new_n712), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n974), .A2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n966), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n970), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n662), .A3(new_n967), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n723), .A2(new_n987), .B1(new_n741), .B2(new_n572), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT111), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n740), .B2(new_n731), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G322), .B2(new_n738), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT48), .Z(new_n1009));
  OAI22_X1  g0809(.A1(new_n979), .A2(new_n746), .B1(new_n991), .B2(new_n735), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n728), .A2(G326), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n254), .B1(new_n791), .B2(G116), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n254), .B1(new_n737), .B2(new_n753), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n731), .A2(new_n269), .B1(new_n741), .B2(new_n203), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n750), .A2(G77), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n724), .A2(G50), .B1(new_n744), .B2(new_n357), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n990), .C1(new_n266), .C2(new_n727), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1017), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n720), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n771), .B1(new_n236), .B2(new_n451), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n665), .A2(new_n223), .A3(new_n254), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n665), .C1(G68), .C2(G77), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n269), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1027), .A2(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n223), .A2(G107), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n777), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n719), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n654), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1026), .A2(new_n712), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1004), .B(new_n1037), .C1(new_n972), .C2(new_n1002), .ZN(G393));
  NAND3_X1  g0838(.A1(new_n954), .A2(new_n655), .A3(new_n960), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n650), .B(new_n654), .C1(new_n953), .C2(new_n959), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n967), .A2(new_n1041), .A3(KEYINPUT115), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(new_n662), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n969), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n967), .A2(new_n1041), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n972), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1039), .A2(new_n1040), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT114), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n777), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n223), .A2(new_n211), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n244), .C2(new_n771), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n744), .A2(G77), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n201), .B2(new_n731), .C1(new_n269), .C2(new_n741), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT112), .Z(new_n1057));
  AOI211_X1 g0857(.A(new_n379), .B(new_n1057), .C1(G143), .C2(new_n728), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n737), .A2(new_n266), .B1(new_n723), .B2(new_n753), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G68), .A2(new_n750), .B1(new_n791), .B2(G87), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n737), .A2(new_n987), .B1(new_n723), .B2(new_n740), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G303), .A2(new_n749), .B1(new_n762), .B2(G294), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n578), .C2(new_n979), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G322), .B2(new_n728), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n379), .C1(new_n746), .C2(new_n735), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1063), .B1(new_n759), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1054), .B1(new_n1070), .B2(new_n720), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n712), .C1(new_n1035), .C2(new_n928), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1050), .A2(new_n1051), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1050), .B2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1048), .B1(new_n1073), .B2(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n684), .A2(new_n644), .A3(new_n785), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n782), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n837), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n869), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n867), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n869), .B1(new_n836), .B2(new_n837), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n868), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n884), .A2(new_n649), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n704), .A2(new_n707), .A3(G330), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n707), .B1(new_n704), .B2(G330), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n878), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(new_n1080), .C1(new_n1081), .C2(new_n868), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1049), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n867), .A2(new_n858), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n859), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n717), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT54), .B(G143), .Z(new_n1094));
  AOI22_X1  g0894(.A1(G128), .A2(new_n738), .B1(new_n762), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n724), .A2(G132), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G125), .B2(new_n728), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n749), .A2(G137), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n750), .A2(G150), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1100), .A2(KEYINPUT53), .B1(new_n753), .B2(new_n979), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(KEYINPUT53), .B2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n254), .B1(new_n747), .B2(new_n201), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT118), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1098), .A2(new_n1099), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1055), .B1(new_n211), .B2(new_n741), .C1(new_n746), .C2(new_n737), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G116), .B2(new_n724), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G87), .A2(new_n750), .B1(new_n791), .B2(G68), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n254), .B1(new_n728), .B2(G294), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n731), .A2(new_n469), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n720), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n806), .A2(new_n269), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1093), .A2(new_n712), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n904), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n685), .B1(new_n811), .B2(new_n671), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT98), .B1(new_n1117), .B2(new_n439), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n613), .B(new_n1116), .C1(new_n1118), .C2(new_n820), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n892), .A2(G330), .A3(new_n812), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n834), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1076), .A2(new_n782), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n812), .B1(new_n832), .B2(new_n833), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n706), .B2(new_n708), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n1123), .A4(new_n1122), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT116), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n812), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1083), .B1(new_n1131), .B2(new_n834), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1132), .B2(new_n829), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n837), .B1(new_n709), .B2(new_n812), .ZN(new_n1134));
  OAI211_X1 g0934(.A(KEYINPUT116), .B(new_n836), .C1(new_n1134), .C2(new_n1083), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1119), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n867), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1079), .B1(new_n829), .B2(new_n834), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1092), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1083), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1088), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1119), .A2(new_n1088), .A3(new_n1084), .A4(new_n1136), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n662), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1089), .B(new_n1115), .C1(new_n1143), .C2(new_n1145), .ZN(G378));
  NOR2_X1   g0946(.A1(new_n290), .A2(new_n291), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n847), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n301), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n611), .A2(new_n282), .A3(new_n1148), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n903), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n891), .A2(new_n894), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT119), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1152), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1153), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1158), .A2(G330), .A3(new_n900), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1157), .A2(new_n1166), .A3(KEYINPUT120), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT120), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n903), .A2(new_n1168), .A3(new_n1156), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1167), .A2(new_n871), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n871), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1049), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n806), .A2(new_n201), .ZN(new_n1173));
  INV_X1    g0973(.A(G125), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n979), .A2(new_n266), .B1(new_n1174), .B2(new_n737), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n724), .A2(G128), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n741), .B2(new_n796), .C1(new_n800), .C2(new_n731), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n750), .C2(new_n1094), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n304), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G41), .B(new_n1181), .C1(G124), .C2(new_n728), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n1179), .B2(new_n1178), .C1(new_n753), .C2(new_n747), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1021), .B1(new_n727), .B2(new_n746), .C1(new_n578), .C2(new_n737), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1184), .A2(new_n254), .A3(new_n980), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n358), .A2(new_n741), .B1(new_n211), .B2(new_n731), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G41), .B(new_n1186), .C1(G58), .C2(new_n791), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(new_n469), .C2(new_n723), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1183), .B(new_n1189), .C1(G50), .C2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n716), .B1(new_n1191), .B2(new_n720), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1173), .B(new_n1192), .C1(new_n1165), .C2(new_n718), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1172), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1165), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT120), .B1(new_n903), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1156), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n895), .B2(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1169), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n871), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1167), .A2(new_n871), .A3(new_n1169), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1202), .A2(new_n1203), .B1(new_n1144), .B2(new_n1119), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n662), .B1(new_n1204), .B2(KEYINPUT57), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1129), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1119), .B1(new_n1142), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(KEYINPUT57), .B(new_n1207), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1195), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT121), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n663), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1194), .B1(new_n1215), .B2(new_n1208), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1212), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(KEYINPUT122), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1119), .B2(new_n1136), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n614), .B(new_n904), .C1(new_n821), .C2(new_n822), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1206), .A2(new_n1221), .A3(KEYINPUT122), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n949), .A3(new_n1137), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT123), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n834), .A2(new_n717), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G283), .A2(new_n724), .B1(new_n728), .B2(G303), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n738), .A2(G294), .B1(new_n744), .B2(new_n357), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n469), .C2(new_n741), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n379), .B1(new_n747), .B2(new_n209), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n578), .B2(new_n731), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1229), .B(new_n1232), .C1(G97), .C2(new_n750), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n749), .A2(new_n1094), .B1(new_n728), .B2(G128), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n254), .C1(new_n266), .C2(new_n741), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G137), .A2(new_n724), .B1(new_n791), .B2(G58), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n753), .B2(new_n735), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n737), .A2(new_n800), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n979), .A2(new_n201), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n720), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n806), .A2(new_n203), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1226), .A2(new_n712), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1206), .B2(new_n972), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1225), .A2(new_n1245), .ZN(G381));
  NOR2_X1   g1046(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1089), .A2(new_n1115), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1212), .A2(new_n1217), .A3(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1048), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n974), .A2(new_n1000), .A3(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT125), .ZN(new_n1255));
  OR4_X1    g1055(.A1(G381), .A2(new_n1250), .A3(new_n1253), .A4(new_n1255), .ZN(G407));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  XOR2_X1   g1057(.A(G393), .B(G396), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1252), .B1(new_n974), .B2(new_n1000), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1000), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(G390), .A2(new_n973), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G390), .B1(new_n973), .B2(new_n1261), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1264), .A3(new_n1258), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1206), .A2(new_n1221), .A3(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n662), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT60), .B1(new_n1206), .B2(new_n1221), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1223), .B2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT126), .B(G384), .C1(new_n1271), .C2(new_n1244), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1119), .A2(new_n1136), .A3(new_n1219), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT122), .B1(new_n1206), .B2(new_n1221), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1270), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1269), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1277), .A2(new_n1245), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G2897), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1272), .A2(new_n1280), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1216), .A2(new_n1249), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1282), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n949), .B(new_n1207), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1172), .A3(new_n1193), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1290), .B2(G378), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1285), .A2(new_n1286), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1210), .B2(G378), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(KEYINPUT62), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1289), .A2(new_n1172), .A3(new_n1193), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1282), .B1(new_n1298), .B2(new_n1249), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1295), .B(new_n1299), .C1(new_n1249), .C2(new_n1216), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1267), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1267), .A2(KEYINPUT61), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1300), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT63), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1283), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1295), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1284), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1210), .A2(G378), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1299), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1308), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1305), .B(new_n1307), .C1(new_n1314), .C2(new_n1306), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(new_n1315), .ZN(G405));
  AND3_X1   g1116(.A1(new_n1250), .A2(new_n1266), .A3(new_n1312), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1266), .B1(new_n1250), .B2(new_n1312), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1295), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1295), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1211), .B(new_n1194), .C1(new_n1215), .C2(new_n1208), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n662), .A3(new_n1208), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT121), .B1(new_n1323), .B2(new_n1195), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1321), .A2(new_n1324), .A3(G378), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1267), .B1(new_n1325), .B2(new_n1287), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1250), .A2(new_n1266), .A3(new_n1312), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1320), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1319), .A2(new_n1328), .ZN(G402));
endmodule


