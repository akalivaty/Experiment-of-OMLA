//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G221), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT12), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT11), .B1(new_n195), .B2(G134), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G137), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n201), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n200), .A4(new_n202), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n202), .A3(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n212), .B(G146), .C1(new_n213), .C2(KEYINPUT1), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n215), .A3(G143), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n214), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT69), .B1(new_n214), .B2(new_n216), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(G143), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n217), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G107), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G104), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT80), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G107), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G104), .B2(new_n224), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT80), .B(G104), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n237), .B(G101), .C1(new_n238), .C2(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G143), .B(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n219), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n214), .A3(new_n216), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n234), .A3(new_n239), .ZN(new_n245));
  AOI221_X4 g059(.A(new_n194), .B1(new_n209), .B2(new_n211), .C1(new_n241), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n228), .A2(KEYINPUT80), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n226), .A2(G104), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n224), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n235), .A3(G104), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G107), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n249), .A2(new_n253), .A3(G101), .ZN(new_n254));
  AOI21_X1  g068(.A(G107), .B1(new_n247), .B2(new_n248), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n255), .A2(new_n231), .A3(new_n236), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n218), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n214), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n243), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n245), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n211), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT12), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n246), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n242), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT0), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n213), .A3(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT0), .B2(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n267), .B1(new_n273), .B2(new_n242), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n251), .B(new_n252), .C1(new_n238), .C2(new_n224), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT81), .A2(G101), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n234), .A2(KEYINPUT4), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT4), .B(new_n278), .C1(new_n249), .C2(new_n253), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n275), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n203), .A2(new_n208), .B1(G131), .B2(new_n210), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n260), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT10), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n245), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(G110), .ZN(new_n292));
  INV_X1    g106(.A(G140), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n266), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n286), .A3(new_n284), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n264), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n298), .B2(new_n287), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n193), .B(new_n189), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n294), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n249), .A2(new_n253), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(new_n231), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n278), .B1(new_n249), .B2(new_n253), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n280), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n217), .A2(new_n218), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n285), .B1(new_n310), .B2(new_n243), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n309), .A2(new_n275), .B1(new_n257), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n283), .B1(new_n312), .B2(new_n286), .ZN(new_n313));
  INV_X1    g127(.A(new_n287), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n303), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n287), .B(new_n294), .C1(new_n246), .C2(new_n265), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n317), .A2(KEYINPUT82), .A3(new_n193), .A4(new_n189), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n303), .B1(new_n266), .B2(new_n314), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n287), .A3(new_n294), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n189), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G469), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n192), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G237), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n288), .A3(G214), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n212), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(new_n288), .A3(G143), .A4(G214), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT18), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n200), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n293), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT86), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n215), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n337), .A2(G146), .ZN(new_n342));
  OAI221_X1 g156(.A(new_n331), .B1(new_n333), .B2(new_n330), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT19), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n337), .A2(KEYINPUT19), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n328), .A2(new_n200), .A3(new_n329), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n351));
  OR3_X1    g165(.A1(new_n335), .A2(KEYINPUT16), .A3(G140), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G146), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n343), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(G113), .B(G122), .Z(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT87), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(G104), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n352), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n215), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(new_n215), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT17), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n333), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n333), .A2(new_n367), .A3(new_n349), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(KEYINPUT88), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n358), .B(new_n343), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G475), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n189), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(KEYINPUT88), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n369), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n366), .C1(new_n370), .C2(new_n369), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n358), .B1(new_n382), .B2(new_n343), .ZN(new_n383));
  INV_X1    g197(.A(new_n374), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n189), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G475), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n375), .A2(KEYINPUT20), .A3(new_n376), .A4(new_n189), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G122), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G116), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n235), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n212), .A2(G128), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n213), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  OAI21_X1  g214(.A(G134), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n398), .A2(new_n395), .A3(new_n201), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n394), .A2(new_n401), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT90), .B1(new_n390), .B2(KEYINPUT14), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n390), .A2(KEYINPUT14), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n389), .A4(G122), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n407), .A2(new_n392), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G107), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n393), .A2(new_n235), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n201), .B1(new_n398), .B2(new_n395), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n413), .B(new_n414), .C1(new_n402), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n188), .A2(G217), .A3(new_n288), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n418), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n406), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n189), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n423), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G234), .A2(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(G952), .A3(new_n288), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT21), .B(G898), .Z(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(G902), .A3(G953), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n388), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G214), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(G110), .B(G122), .Z(new_n439));
  XOR2_X1   g253(.A(KEYINPUT2), .B(G113), .Z(new_n440));
  XNOR2_X1  g254(.A(G116), .B(G119), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(KEYINPUT2), .A2(G113), .ZN(new_n443));
  INV_X1    g257(.A(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n389), .A2(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT2), .A2(G113), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(KEYINPUT70), .A3(new_n441), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n307), .B1(new_n254), .B2(new_n304), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(new_n280), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT83), .B1(new_n445), .B2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n444), .A4(G116), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(G113), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n240), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n439), .B1(new_n454), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n440), .A2(new_n441), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n279), .B2(new_n281), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n257), .A2(new_n455), .A3(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(new_n439), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n274), .A2(G125), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n258), .A2(new_n335), .A3(new_n243), .A4(new_n259), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n288), .A2(G224), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT84), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n474), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n439), .C1(new_n454), .C2(new_n463), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(KEYINPUT7), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n472), .B2(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n439), .B(KEYINPUT8), .Z(new_n486));
  AND2_X1   g300(.A1(new_n462), .A2(new_n240), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n463), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n472), .A2(new_n473), .A3(new_n482), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n470), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n189), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n480), .A2(new_n490), .A3(new_n189), .A4(new_n492), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n438), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n325), .A2(new_n436), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n283), .B2(new_n274), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n195), .A2(G134), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n200), .B1(new_n500), .B2(new_n202), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT68), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n209), .A2(new_n260), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n264), .A2(KEYINPUT67), .A3(new_n275), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n264), .A2(new_n275), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT30), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n466), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n452), .A3(new_n503), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n326), .A2(new_n288), .A3(G210), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT27), .Z(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT26), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n231), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT31), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n512), .A2(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n505), .A2(new_n466), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n518), .ZN(new_n525));
  INV_X1    g339(.A(new_n512), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n505), .A2(new_n506), .B1(new_n509), .B2(KEYINPUT30), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n466), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n517), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n523), .A3(new_n517), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n528), .C2(new_n517), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n509), .A2(new_n452), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n520), .B2(new_n521), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT29), .A3(new_n517), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n541), .A2(KEYINPUT71), .A3(KEYINPUT29), .A4(new_n517), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n539), .A2(new_n544), .A3(new_n189), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G472), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n536), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n353), .B1(G146), .B2(new_n337), .ZN(new_n550));
  XNOR2_X1  g364(.A(G119), .B(G128), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT23), .B1(new_n213), .B2(G119), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT73), .B1(new_n213), .B2(G119), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  OR3_X1    g376(.A1(new_n561), .A2(new_n562), .A3(G110), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n550), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n566));
  OAI21_X1  g380(.A(G110), .B1(new_n561), .B2(new_n562), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n363), .A2(new_n566), .A3(new_n365), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT76), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n195), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(G137), .A3(new_n575), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n363), .A2(new_n365), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(KEYINPUT75), .A3(new_n566), .A4(new_n567), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n568), .A2(new_n569), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n581), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n565), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n549), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n586), .B2(new_n565), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n564), .B(new_n581), .C1(new_n584), .C2(new_n585), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n189), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n595));
  INV_X1    g409(.A(G217), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(G234), .B2(new_n189), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n582), .A2(new_n588), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n497), .A2(new_n548), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n531), .A2(new_n189), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(G472), .B1(new_n532), .B2(new_n531), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n603), .A3(new_n325), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n494), .A2(new_n495), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT92), .B1(new_n609), .B2(new_n437), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n611), .B(new_n438), .C1(new_n494), .C2(new_n495), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n419), .A2(KEYINPUT33), .A3(new_n421), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT33), .B1(new_n419), .B2(new_n421), .ZN(new_n615));
  OAI21_X1  g429(.A(G478), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n422), .A2(new_n424), .A3(new_n189), .ZN(new_n617));
  NAND2_X1  g431(.A1(G478), .A2(G902), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT93), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT93), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n616), .A2(new_n621), .A3(new_n617), .A4(new_n618), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n388), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n613), .A2(new_n434), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n608), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND4_X1  g442(.A1(new_n379), .A2(new_n429), .A3(new_n386), .A4(new_n387), .ZN(new_n629));
  OR3_X1    g443(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n435), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n629), .B2(new_n435), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n613), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n608), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT35), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G107), .ZN(G9));
  NAND2_X1  g450(.A1(new_n606), .A2(G472), .ZN(new_n637));
  INV_X1    g451(.A(new_n572), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n600), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n598), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n637), .A2(new_n533), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n607), .A2(KEYINPUT96), .A3(new_n643), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n497), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT97), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AND2_X1   g465(.A1(new_n325), .A2(new_n643), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n288), .A2(G900), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n430), .A2(G902), .ZN(new_n655));
  OR3_X1    g469(.A1(new_n654), .A2(KEYINPUT98), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n431), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n629), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n652), .A2(new_n548), .A3(new_n613), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XNOR2_X1  g476(.A(new_n658), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT39), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n325), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n643), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n609), .B(KEYINPUT38), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n429), .A3(new_n388), .A4(new_n437), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n528), .A2(new_n518), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n518), .A2(new_n512), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n189), .B1(new_n675), .B2(new_n540), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n535), .A2(new_n536), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n670), .A2(new_n682), .A3(new_n673), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n212), .ZN(G45));
  NOR2_X1   g499(.A1(new_n623), .A2(new_n659), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n652), .A2(new_n548), .A3(new_n613), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(new_n625), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT32), .B1(new_n531), .B2(new_n532), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n602), .B1(new_n692), .B2(new_n547), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n189), .B1(new_n296), .B2(new_n299), .ZN(new_n694));
  AOI221_X4 g508(.A(new_n192), .B1(G469), .B2(new_n694), .C1(new_n302), .C2(new_n318), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND3_X1  g512(.A1(new_n548), .A2(new_n603), .A3(new_n695), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n632), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n389), .ZN(G18));
  AND2_X1   g515(.A1(new_n643), .A2(new_n436), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n609), .A2(new_n437), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n611), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n496), .A2(KEYINPUT92), .ZN(new_n705));
  AND4_X1   g519(.A1(KEYINPUT103), .A2(new_n695), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT103), .B1(new_n613), .B2(new_n695), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n548), .B(new_n702), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NAND2_X1  g523(.A1(new_n388), .A2(new_n429), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n610), .A2(new_n612), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n434), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT104), .B(G472), .Z(new_n713));
  OAI211_X1 g527(.A(new_n519), .B(new_n530), .C1(new_n517), .C2(new_n541), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n606), .A2(new_n713), .B1(new_n532), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n603), .A3(new_n695), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT105), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND3_X1  g533(.A1(new_n715), .A2(new_n686), .A3(new_n643), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n695), .A2(new_n704), .A3(new_n705), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n613), .A2(KEYINPUT103), .A3(new_n695), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n335), .ZN(G27));
  NOR2_X1   g540(.A1(new_n192), .A2(new_n438), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n494), .A2(new_n495), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n319), .A2(new_n324), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n319), .A2(KEYINPUT106), .A3(new_n324), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n548), .A3(new_n603), .A4(new_n686), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT107), .A3(KEYINPUT42), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n736));
  NAND4_X1  g550(.A1(new_n693), .A2(new_n686), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n200), .ZN(G33));
  NAND4_X1  g553(.A1(new_n733), .A2(new_n548), .A3(new_n603), .A4(new_n660), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  XNOR2_X1  g555(.A(new_n322), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(G469), .C1(new_n742), .C2(G902), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n319), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n191), .A3(new_n665), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n620), .A2(new_n622), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n388), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT43), .ZN(new_n752));
  INV_X1    g566(.A(new_n607), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n643), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n609), .A2(new_n438), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n753), .A4(new_n643), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND3_X1  g574(.A1(new_n692), .A2(new_n547), .A3(new_n602), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n686), .A2(new_n757), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n748), .A2(new_n191), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n748), .A2(new_n768), .A3(new_n191), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n764), .A2(new_n765), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT99), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n678), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n694), .A2(G469), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n319), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n431), .A3(new_n728), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n773), .A2(new_n603), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n624), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n288), .A2(G952), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n693), .A2(new_n752), .A3(new_n776), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n778), .B(new_n782), .C1(new_n781), .C2(new_n780), .ZN(new_n783));
  INV_X1    g597(.A(new_n388), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n784), .A3(new_n750), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n716), .ZN(new_n788));
  INV_X1    g602(.A(new_n431), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n671), .A2(new_n437), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n752), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n791), .B(new_n793), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n752), .A2(new_n789), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n715), .A2(new_n603), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n767), .A2(new_n769), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n775), .A2(new_n191), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n757), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n752), .A2(new_n643), .A3(new_n715), .A4(new_n776), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n787), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT51), .B1(new_n801), .B2(KEYINPUT117), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n783), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n715), .A2(new_n643), .A3(new_n686), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n706), .B2(new_n707), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n598), .A2(new_n642), .A3(new_n658), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n731), .B2(new_n732), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n191), .A3(new_n678), .A4(new_n711), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n661), .A3(new_n687), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT109), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n548), .A2(new_n652), .A3(new_n613), .A4(new_n660), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n725), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n812), .A2(new_n687), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n699), .A2(new_n625), .B1(new_n712), .B2(new_n716), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n548), .A2(new_n702), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n723), .B2(new_n724), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n826), .A3(new_n700), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n735), .A2(new_n737), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT112), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  INV_X1    g644(.A(new_n632), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n693), .A3(new_n695), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n696), .A2(new_n708), .A3(new_n832), .A4(new_n717), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n833), .B2(new_n738), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n435), .B(new_n703), .C1(new_n623), .C2(new_n629), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n603), .A3(new_n325), .A4(new_n607), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n648), .A2(new_n604), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n808), .A2(new_n733), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n388), .A2(new_n429), .A3(new_n659), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n652), .A2(new_n548), .A3(new_n757), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n839), .A2(new_n840), .A3(new_n844), .A4(new_n740), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n648), .A2(new_n604), .A3(new_n838), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n740), .A3(new_n843), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT111), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n836), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n823), .A2(new_n835), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n814), .A2(new_n819), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n833), .A2(new_n738), .A3(new_n846), .A4(new_n847), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n814), .A2(new_n819), .A3(KEYINPUT52), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n836), .ZN(new_n859));
  XOR2_X1   g673(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n823), .A2(new_n835), .A3(new_n849), .A4(KEYINPUT113), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n852), .A2(new_n859), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n823), .A2(new_n836), .A3(new_n856), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n807), .A2(new_n867), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n796), .B(new_n795), .C1(new_n723), .C2(new_n724), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n868), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n775), .B(KEYINPUT49), .Z(new_n871));
  NOR4_X1   g685(.A1(new_n671), .A2(new_n602), .A3(new_n388), .A4(new_n750), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n773), .A2(new_n727), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(G75));
  NAND3_X1  g688(.A1(new_n852), .A2(new_n859), .A3(new_n862), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(G210), .A3(G902), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n471), .A2(new_n479), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n477), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n288), .A2(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n860), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n863), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(new_n744), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n744), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n317), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n875), .A2(G469), .A3(G902), .A4(new_n742), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n891), .B2(new_n892), .ZN(G54));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT119), .B1(new_n894), .B2(new_n376), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n894), .A2(new_n376), .A3(KEYINPUT119), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n875), .A2(G902), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n375), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n883), .ZN(G60));
  NOR2_X1   g715(.A1(new_n614), .A2(new_n615), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n618), .B(KEYINPUT59), .Z(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n886), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  INV_X1    g721(.A(new_n883), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n905), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n885), .B2(new_n863), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT120), .B1(new_n911), .B2(new_n883), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n863), .B2(new_n866), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n913), .B2(new_n902), .ZN(new_n914));
  INV_X1    g728(.A(new_n904), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n867), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n903), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n909), .A2(new_n912), .B1(new_n914), .B2(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n875), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n599), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n875), .A2(new_n641), .A3(new_n921), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n908), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G66));
  NAND2_X1  g742(.A1(new_n432), .A2(G224), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G953), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n833), .A2(new_n846), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n878), .B1(G898), .B2(new_n288), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G69));
  INV_X1    g748(.A(G227), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n653), .B1(new_n935), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT124), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n347), .B(KEYINPUT122), .Z(new_n939));
  XOR2_X1   g753(.A(new_n527), .B(new_n939), .Z(new_n940));
  AND2_X1   g754(.A1(new_n759), .A2(new_n770), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n602), .B(new_n749), .C1(new_n692), .C2(new_n547), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n738), .B1(new_n942), .B2(new_n711), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n816), .A2(new_n687), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n941), .A2(new_n943), .A3(new_n740), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n288), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT125), .B1(new_n946), .B2(new_n654), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n948), .B(new_n653), .C1(new_n945), .C2(new_n288), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n940), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n940), .C1(new_n947), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n681), .A2(new_n944), .A3(new_n683), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n681), .A2(new_n944), .A3(KEYINPUT62), .A4(new_n683), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n623), .A2(new_n629), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n693), .A2(new_n666), .A3(new_n757), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n961), .A3(new_n941), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n940), .B1(new_n962), .B2(new_n288), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n938), .B1(new_n954), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT123), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n937), .B(new_n965), .C1(new_n966), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  INV_X1    g784(.A(new_n931), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n883), .B1(new_n972), .B2(new_n674), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n945), .B2(new_n971), .ZN(new_n974));
  INV_X1    g788(.A(new_n675), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n511), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n674), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n511), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n864), .A2(new_n977), .A3(new_n865), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n970), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n973), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT127), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n973), .A2(new_n985), .A3(new_n982), .A4(new_n976), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G57));
endmodule


