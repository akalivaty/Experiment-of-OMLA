//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n189), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n194), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT66), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n195), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT64), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n210), .A2(G134), .ZN(new_n215));
  OAI211_X1 g029(.A(G131), .B(new_n211), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n213), .B2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(G137), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n224), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n228), .B(KEYINPUT1), .C1(new_n229), .C2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n227), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n223), .B1(new_n226), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  OR2_X1    g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n229), .A2(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n232), .A2(G143), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n237), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n229), .A2(G146), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n233), .A2(new_n242), .A3(KEYINPUT0), .A4(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n222), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n209), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n235), .A2(new_n226), .ZN(new_n250));
  INV_X1    g064(.A(new_n223), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT66), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n191), .B2(new_n193), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n255), .A2(new_n195), .B1(new_n196), .B2(new_n203), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n246), .A2(new_n222), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n243), .A3(new_n241), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n248), .A2(new_n249), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT28), .B1(new_n248), .B2(new_n249), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n188), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n256), .B1(new_n252), .B2(new_n258), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(KEYINPUT70), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n248), .A2(new_n249), .A3(new_n259), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n259), .A2(new_n268), .A3(new_n263), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n259), .B2(new_n263), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G237), .A2(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G210), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT27), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G101), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n277), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n259), .A2(new_n282), .A3(new_n277), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(KEYINPUT30), .C1(new_n236), .C2(new_n247), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n285), .A2(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(KEYINPUT30), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n252), .A2(new_n258), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n256), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n279), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n259), .A2(new_n282), .A3(new_n277), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n282), .B1(new_n259), .B2(new_n277), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n286), .A2(new_n289), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n209), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n272), .A2(new_n278), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n187), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n270), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n259), .A2(new_n268), .A3(new_n263), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT71), .B1(new_n265), .B2(new_n266), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n277), .B1(new_n306), .B2(new_n267), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT31), .B1(new_n294), .B2(new_n296), .ZN(new_n308));
  NOR4_X1   g122(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(new_n279), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(KEYINPUT73), .B(new_n299), .C1(new_n307), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n301), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n272), .A2(new_n278), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n291), .A2(new_n297), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n300), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n262), .A2(new_n277), .A3(new_n267), .A4(new_n271), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n296), .A2(new_n259), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n318), .B2(new_n278), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n248), .A2(new_n259), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT28), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n271), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G902), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(KEYINPUT32), .A2(new_n316), .B1(new_n327), .B2(G472), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n313), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT16), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n332), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G146), .ZN(new_n336));
  XNOR2_X1  g150(.A(G125), .B(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n232), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n190), .B2(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n342));
  INV_X1    g156(.A(G110), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n340), .B(new_n344), .C1(new_n190), .C2(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n190), .A2(G128), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G119), .B(G128), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT24), .B(G110), .Z(new_n349));
  OAI22_X1  g163(.A1(new_n347), .A2(KEYINPUT76), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n339), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n334), .A2(new_n335), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n232), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n336), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n356), .A2(G110), .B1(new_n348), .B2(new_n349), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n355), .B2(new_n357), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  INV_X1    g176(.A(G953), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(G221), .A3(G234), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n356), .A2(G110), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n349), .A2(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n336), .ZN(new_n371));
  AOI21_X1  g185(.A(G146), .B1(new_n334), .B2(new_n335), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT75), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n352), .A3(new_n365), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n377), .A3(new_n325), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n367), .A2(new_n377), .A3(KEYINPUT25), .A4(new_n325), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G217), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G234), .B2(new_n325), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n367), .A2(new_n377), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n384), .A2(G902), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n384), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n380), .B2(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(new_n389), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT77), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n329), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G210), .B1(G237), .B2(G902), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT87), .Z(new_n399));
  OAI21_X1  g213(.A(KEYINPUT5), .B1(new_n253), .B2(new_n254), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n403), .A2(new_n190), .A3(KEYINPUT84), .A4(G116), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n402), .A2(G113), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n400), .A2(new_n405), .B1(new_n196), .B2(new_n203), .ZN(new_n406));
  INV_X1    g220(.A(G104), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G104), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT3), .B1(new_n407), .B2(G107), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(KEYINPUT3), .C1(new_n407), .C2(G107), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT80), .B(G101), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n407), .A2(KEYINPUT81), .A3(G107), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n410), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n416), .A2(new_n417), .B1(G101), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G101), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT4), .B1(new_n416), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n409), .A2(G104), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n407), .A2(G107), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n414), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n430));
  INV_X1    g244(.A(new_n415), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n429), .B(new_n417), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G101), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n209), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n423), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n423), .B(new_n440), .C1(new_n434), .C2(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n413), .A2(new_n415), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n424), .B1(new_n445), .B2(new_n429), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n436), .A2(new_n446), .B1(new_n204), .B2(new_n208), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n432), .B(KEYINPUT4), .C1(new_n424), .C2(new_n416), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n422), .B2(new_n406), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n440), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n235), .A2(new_n332), .A3(new_n226), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n244), .A2(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G224), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n444), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n440), .B(KEYINPUT8), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n403), .B1(new_n206), .B2(new_n207), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n402), .A2(G113), .A3(new_n404), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n204), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n462), .B2(new_n422), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n421), .A2(G101), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n432), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(G113), .A3(new_n402), .A4(new_n404), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n204), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n458), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n406), .A2(new_n465), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n204), .A2(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n422), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT85), .A4(new_n459), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n453), .A2(new_n475), .A3(new_n455), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n449), .B2(new_n440), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n452), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n479), .A2(new_n480), .B1(new_n475), .B2(new_n455), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n325), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n399), .B1(new_n457), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n444), .A2(new_n450), .A3(new_n456), .ZN(new_n486));
  INV_X1    g300(.A(new_n399), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n325), .A3(new_n487), .A4(new_n482), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT88), .B(new_n399), .C1(new_n457), .C2(new_n483), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT9), .B(G234), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(new_n383), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n496));
  INV_X1    g310(.A(G128), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(G143), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n229), .A2(KEYINPUT95), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(KEYINPUT13), .A3(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(G143), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G134), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n192), .B2(G122), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT94), .A3(G116), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n192), .A2(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G107), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n508), .A2(new_n510), .B1(new_n192), .B2(G122), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n409), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n500), .A2(new_n213), .A3(new_n504), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n409), .B1(new_n511), .B2(new_n512), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(KEYINPUT14), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n515), .B1(KEYINPUT14), .B2(new_n409), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n500), .A2(new_n213), .A3(new_n504), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n213), .B1(new_n500), .B2(new_n504), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n519), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n520), .B1(new_n519), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n495), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n500), .A2(new_n501), .B1(new_n497), .B2(G143), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n213), .B1(new_n531), .B2(new_n503), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n511), .A2(new_n409), .A3(new_n512), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n518), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n521), .A2(new_n522), .ZN(new_n536));
  OAI22_X1  g350(.A1(new_n532), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT96), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n519), .A2(new_n527), .A3(new_n520), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n494), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n530), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n325), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n541), .B(new_n325), .C1(KEYINPUT15), .C2(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G237), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n363), .A3(G214), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n229), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n273), .A2(G143), .A3(G214), .ZN(new_n552));
  NAND2_X1  g366(.A1(KEYINPUT18), .A2(G131), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n551), .A2(KEYINPUT89), .A3(new_n552), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n331), .A2(new_n333), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G146), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n338), .ZN(new_n560));
  INV_X1    g374(.A(new_n553), .ZN(new_n561));
  INV_X1    g375(.A(new_n552), .ZN(new_n562));
  AOI21_X1  g376(.A(G143), .B1(new_n273), .B2(G214), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n556), .A2(new_n557), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT90), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n551), .A2(new_n552), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n561), .B1(new_n559), .B2(new_n338), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n569), .A2(KEYINPUT90), .A3(new_n557), .A4(new_n556), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G113), .B(G122), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n407), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(KEYINPUT17), .A3(G131), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n574), .A2(new_n354), .A3(new_n336), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(G131), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n551), .A2(new_n220), .A3(new_n552), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n567), .A2(new_n570), .B1(new_n579), .B2(new_n575), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT92), .A3(new_n573), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n578), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n337), .B(KEYINPUT19), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n371), .B1(new_n587), .B2(new_n232), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n567), .A2(new_n570), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n573), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n586), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n571), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT91), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n583), .A2(new_n585), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G475), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT20), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT92), .B1(new_n584), .B2(new_n573), .ZN(new_n599));
  AND4_X1   g413(.A1(KEYINPUT92), .A2(new_n571), .A3(new_n573), .A4(new_n580), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n571), .A2(new_n590), .A3(new_n592), .ZN(new_n601));
  INV_X1    g415(.A(new_n573), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n589), .A2(new_n590), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n599), .A2(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n596), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n584), .A2(new_n573), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n583), .B2(new_n585), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT93), .B1(new_n610), .B2(G902), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n584), .A2(new_n573), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(new_n600), .B2(new_n599), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n325), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n615), .A3(G475), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n548), .A2(new_n608), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G221), .B1(new_n493), .B2(G902), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT78), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n244), .B1(new_n446), .B2(new_n436), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n448), .ZN(new_n621));
  INV_X1    g435(.A(new_n257), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n422), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n497), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n226), .B1(new_n624), .B2(new_n224), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n432), .A2(new_n625), .A3(new_n464), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n626), .B1(new_n422), .B2(new_n250), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n630), .A2(KEYINPUT12), .A3(new_n257), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT12), .B1(new_n630), .B2(new_n257), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(G110), .B(G140), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n363), .A2(G227), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n629), .A2(KEYINPUT82), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n621), .A2(new_n623), .A3(new_n628), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n257), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT82), .B1(new_n629), .B2(new_n638), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT83), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n637), .B(KEYINPUT83), .C1(new_n642), .C2(new_n643), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(G469), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G469), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n325), .ZN(new_n650));
  INV_X1    g464(.A(new_n629), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n620), .A2(new_n448), .B1(new_n626), .B2(new_n627), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n622), .B1(new_n652), .B2(new_n623), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n636), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n629), .B(new_n638), .C1(new_n631), .C2(new_n632), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n650), .B1(new_n656), .B2(new_n649), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n619), .B1(new_n648), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(G214), .B1(G237), .B2(G902), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(G234), .A2(G237), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(G902), .A3(G953), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT21), .B(G898), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n363), .A2(G952), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(G234), .B2(G237), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n660), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n492), .A2(new_n617), .A3(new_n658), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n397), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n417), .ZN(G3));
  AND2_X1   g487(.A1(new_n301), .A2(new_n311), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n396), .A3(new_n658), .A4(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n660), .B1(new_n484), .B2(new_n488), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n665), .A2(new_n668), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n608), .A2(new_n616), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT33), .ZN(new_n683));
  INV_X1    g497(.A(new_n540), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n494), .B1(new_n538), .B2(new_n539), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n541), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n530), .A2(KEYINPUT33), .A3(new_n540), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n530), .A2(KEYINPUT100), .A3(new_n540), .A4(KEYINPUT33), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n688), .A2(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n543), .A2(G902), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n694), .A2(new_n695), .B1(new_n543), .B2(new_n542), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n680), .A2(new_n682), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n677), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT34), .B(G104), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G6));
  INV_X1    g514(.A(new_n680), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n606), .B1(new_n605), .B2(new_n596), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT101), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n547), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n616), .A2(KEYINPUT102), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n611), .A2(new_n615), .A3(new_n709), .A4(G475), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n677), .A2(new_n701), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT35), .B(G107), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G9));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n376), .B2(new_n352), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n716), .B(new_n352), .C1(new_n359), .C2(new_n360), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  OAI22_X1  g533(.A1(new_n717), .A2(new_n719), .B1(KEYINPUT36), .B2(new_n366), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n361), .A2(KEYINPUT103), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n718), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n382), .A2(new_n384), .B1(new_n724), .B2(new_n388), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n674), .A2(new_n675), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n670), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT104), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT37), .B(G110), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G12));
  AOI211_X1 g545(.A(new_n619), .B(new_n725), .C1(new_n648), .C2(new_n657), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n329), .A2(new_n732), .A3(new_n678), .ZN(new_n733));
  INV_X1    g547(.A(new_n707), .ZN(new_n734));
  INV_X1    g548(.A(new_n711), .ZN(new_n735));
  INV_X1    g549(.A(G900), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n667), .B1(new_n663), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT105), .B(G128), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G30));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n491), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n682), .A2(new_n548), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n726), .A2(new_n660), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n737), .B(KEYINPUT39), .Z(new_n748));
  NAND2_X1  g562(.A1(new_n658), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT40), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(KEYINPUT40), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n316), .A2(KEYINPUT32), .ZN(new_n752));
  INV_X1    g566(.A(G472), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n325), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n294), .A2(new_n296), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n321), .B2(new_n278), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT107), .Z(new_n758));
  NAND3_X1  g572(.A1(new_n313), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n747), .A2(new_n750), .A3(new_n751), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G143), .ZN(G45));
  NAND2_X1  g575(.A1(new_n692), .A2(new_n693), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT99), .B1(new_n541), .B2(new_n683), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n687), .B(KEYINPUT33), .C1(new_n530), .C2(new_n540), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n762), .B(new_n695), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n542), .A2(new_n543), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(new_n681), .A3(new_n738), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n329), .A3(new_n678), .A4(new_n732), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G146), .ZN(G48));
  AOI21_X1  g584(.A(new_n395), .B1(new_n313), .B2(new_n328), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n656), .A2(new_n649), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n656), .A2(new_n649), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n619), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n697), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT41), .B(G113), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G15));
  NAND4_X1  g592(.A1(new_n771), .A2(new_n712), .A3(new_n701), .A4(new_n775), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G116), .ZN(G18));
  INV_X1    g594(.A(new_n775), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n680), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n329), .A3(new_n617), .A4(new_n726), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G119), .ZN(G21));
  NAND2_X1  g598(.A1(new_n271), .A2(new_n322), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n278), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n300), .B1(new_n315), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(G902), .B1(new_n314), .B2(new_n315), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT108), .B1(new_n788), .B2(new_n753), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(G472), .C1(new_n298), .C2(G902), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n392), .A2(new_n393), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n782), .A2(new_n792), .A3(new_n793), .A4(new_n745), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G122), .ZN(G24));
  NAND3_X1  g609(.A1(new_n767), .A2(new_n681), .A3(new_n738), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n775), .A2(new_n678), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n725), .B(new_n787), .C1(new_n789), .C2(new_n791), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G125), .ZN(G27));
  OAI211_X1 g615(.A(new_n637), .B(G469), .C1(new_n642), .C2(new_n643), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n619), .B1(new_n657), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n491), .A2(new_n659), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n771), .A2(new_n804), .A3(new_n768), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n660), .B1(new_n489), .B2(new_n490), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n765), .A2(new_n766), .B1(new_n608), .B2(new_n616), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n738), .A4(new_n803), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n327), .A2(G472), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n312), .B1(new_n298), .B2(new_n300), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n752), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(KEYINPUT42), .A3(new_n793), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT109), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n810), .A2(new_n814), .A3(KEYINPUT109), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n807), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT110), .B(G131), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G33));
  NAND4_X1  g634(.A1(new_n771), .A2(new_n804), .A3(new_n712), .A4(new_n738), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G134), .ZN(G36));
  NAND2_X1  g636(.A1(new_n674), .A2(new_n675), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n726), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n681), .B(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT43), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n696), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n696), .B2(new_n681), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n824), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n808), .B1(new_n831), .B2(KEYINPUT44), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(KEYINPUT44), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n646), .A2(new_n647), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT45), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(G469), .B1(new_n644), .B2(new_n835), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(new_n650), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT46), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n646), .B2(new_n647), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT46), .B(new_n841), .C1(new_n843), .C2(new_n837), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT111), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n772), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT46), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n839), .A2(new_n841), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n846), .A2(KEYINPUT112), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n842), .A2(new_n845), .A3(new_n850), .A4(new_n772), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n619), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n833), .A2(new_n748), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G137), .ZN(G39));
  INV_X1    g668(.A(new_n808), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n329), .A2(new_n855), .A3(new_n796), .A4(new_n396), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT47), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n857), .B(new_n619), .C1(new_n849), .C2(new_n851), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n848), .A2(new_n847), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n851), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n619), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT47), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n856), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(G140), .ZN(G42));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n855), .A2(new_n781), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT117), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n759), .A2(new_n395), .A3(new_n668), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n809), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n668), .B1(new_n829), .B2(new_n830), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n792), .A2(new_n793), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n678), .A3(new_n775), .A4(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n666), .B(KEYINPUT119), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT48), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n813), .A2(new_n793), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n868), .A2(new_n871), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n877), .A3(new_n871), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT48), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n872), .A3(new_n808), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n858), .A2(new_n863), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n773), .A2(new_n774), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n619), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n767), .A2(new_n681), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n869), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n868), .A2(KEYINPUT118), .A3(new_n869), .A4(new_n887), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n744), .A2(new_n659), .A3(new_n781), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n871), .A2(new_n872), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT50), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n871), .A2(new_n895), .A3(KEYINPUT50), .A4(new_n872), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n868), .A2(new_n799), .A3(new_n871), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n894), .A2(new_n900), .A3(KEYINPUT51), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n881), .B1(new_n886), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n861), .A2(new_n862), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n857), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n852), .A2(KEYINPUT47), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n885), .ZN(new_n907));
  INV_X1    g721(.A(new_n882), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT51), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n866), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n886), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n909), .A2(KEYINPUT51), .A3(new_n910), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(KEYINPUT120), .A3(new_n916), .A4(new_n881), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n792), .A2(new_n726), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n809), .A2(new_n678), .A3(new_n738), .A4(new_n775), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n733), .A2(new_n739), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n800), .B(KEYINPUT115), .C1(new_n739), .C2(new_n733), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n681), .A2(new_n547), .A3(new_n678), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n803), .A2(new_n725), .A3(new_n738), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n759), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n769), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT52), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT52), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n769), .A2(new_n926), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n920), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n810), .A2(new_n814), .A3(KEYINPUT109), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n933), .A2(new_n815), .B1(new_n806), .B2(new_n805), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n776), .A2(new_n779), .A3(new_n783), .A4(new_n794), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT53), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT116), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n804), .A2(new_n768), .A3(new_n726), .A4(new_n792), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n821), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n547), .A2(new_n737), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n705), .A2(new_n941), .A3(new_n706), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT114), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n942), .A2(new_n735), .A3(new_n943), .A4(new_n808), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n329), .A2(new_n732), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n735), .A3(new_n808), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(KEYINPUT114), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n670), .B1(new_n397), .B2(new_n727), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n696), .A2(new_n681), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n548), .A2(new_n608), .A3(new_n616), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n492), .A3(new_n951), .A4(new_n669), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n676), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n938), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n821), .A2(new_n939), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n946), .A2(KEYINPUT114), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(new_n329), .A3(new_n732), .A4(new_n944), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n938), .A2(new_n954), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n932), .B(new_n937), .C1(new_n955), .C2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n935), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n948), .A2(new_n818), .A3(new_n961), .A4(new_n954), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n329), .A2(new_n732), .A3(new_n678), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n707), .A2(new_n711), .A3(new_n737), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n963), .A2(new_n964), .B1(new_n799), .B2(new_n798), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT52), .B1(new_n965), .B2(new_n927), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n920), .A2(new_n930), .A3(new_n929), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n936), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT54), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n960), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n948), .A2(new_n954), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n934), .A2(new_n935), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n932), .A3(new_n936), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT53), .B1(new_n962), .B2(new_n968), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT54), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n912), .A2(new_n917), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(G952), .A2(G953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n884), .B(KEYINPUT49), .Z(new_n981));
  NAND3_X1  g795(.A1(new_n793), .A2(new_n862), .A3(new_n659), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n696), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n759), .ZN(new_n984));
  INV_X1    g798(.A(new_n744), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n826), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n980), .A2(new_n986), .ZN(G75));
  NOR2_X1   g801(.A1(new_n363), .A2(G952), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n325), .B1(new_n960), .B2(new_n969), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT56), .B1(new_n990), .B2(new_n399), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n444), .A2(new_n450), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n456), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT55), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n991), .A2(new_n994), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT121), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n991), .A2(KEYINPUT121), .A3(new_n994), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G51));
  NAND2_X1  g814(.A1(new_n960), .A2(new_n969), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT54), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n971), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT122), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1001), .A2(new_n1004), .A3(KEYINPUT54), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n650), .B(KEYINPUT57), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n654), .A2(new_n655), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n990), .A2(new_n836), .A3(new_n838), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .ZN(G54));
  NAND2_X1  g825(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT123), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n990), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n989), .B1(new_n1014), .B2(new_n605), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n605), .B2(new_n1014), .ZN(G60));
  NAND2_X1  g830(.A1(G478), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT59), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n971), .B2(new_n976), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n989), .B1(new_n1019), .B2(new_n694), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1021));
  INV_X1    g835(.A(new_n694), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n1018), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(G63));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT60), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n960), .B2(new_n969), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1027), .A2(new_n387), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n724), .B(KEYINPUT124), .Z(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1028), .A2(new_n989), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT61), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1028), .A2(KEYINPUT61), .A3(new_n989), .A4(new_n1030), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(G66));
  OAI21_X1  g849(.A(G953), .B1(new_n664), .B2(new_n454), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n961), .A2(new_n954), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1036), .B1(new_n1038), .B2(G953), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n992), .B1(G898), .B2(new_n363), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(G69));
  NAND2_X1  g855(.A1(new_n818), .A2(new_n821), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n922), .A2(new_n769), .A3(new_n923), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n852), .A2(new_n748), .A3(new_n877), .A4(new_n924), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n853), .A2(new_n864), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n295), .B(new_n587), .Z(new_n1047));
  NOR2_X1   g861(.A1(new_n1047), .A2(G953), .ZN(new_n1048));
  AOI22_X1  g862(.A1(new_n1046), .A2(new_n1048), .B1(new_n736), .B2(G953), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n853), .A2(new_n864), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n950), .A2(new_n951), .A3(new_n808), .ZN(new_n1051));
  NOR3_X1   g865(.A1(new_n397), .A2(new_n1051), .A3(new_n749), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n760), .A2(new_n922), .A3(new_n769), .A4(new_n923), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT62), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g871(.A(G953), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1047), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1049), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n363), .B1(G227), .B2(G900), .ZN(new_n1061));
  XNOR2_X1  g875(.A(new_n1060), .B(new_n1061), .ZN(G72));
  XNOR2_X1  g876(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1063), .B(new_n754), .Z(new_n1064));
  OAI21_X1  g878(.A(new_n1064), .B1(new_n1046), .B2(new_n1037), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(KEYINPUT126), .ZN(new_n1066));
  INV_X1    g880(.A(KEYINPUT126), .ZN(new_n1067));
  OAI211_X1 g881(.A(new_n1067), .B(new_n1064), .C1(new_n1046), .C2(new_n1037), .ZN(new_n1068));
  NOR2_X1   g882(.A1(new_n318), .A2(new_n277), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g884(.A1(new_n1050), .A2(new_n1057), .A3(new_n1038), .ZN(new_n1071));
  INV_X1    g885(.A(new_n1064), .ZN(new_n1072));
  OAI211_X1 g886(.A(new_n277), .B(new_n318), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n318), .A2(new_n278), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1072), .B1(new_n1074), .B2(new_n755), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n974), .A2(new_n975), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT127), .ZN(new_n1077));
  OR2_X1    g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n988), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g894(.A1(new_n1070), .A2(new_n1073), .A3(new_n1080), .ZN(G57));
endmodule


