

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(KEYINPUT32), .B(KEYINPUT102), .ZN(n753) );
  XNOR2_X1 U554 ( .A(n754), .B(n753), .ZN(n763) );
  AND2_X1 U555 ( .A1(n697), .A2(n696), .ZN(n698) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U557 ( .A(n726), .B(n725), .ZN(n732) );
  XNOR2_X1 U558 ( .A(n744), .B(KEYINPUT100), .ZN(n755) );
  NOR2_X2 U559 ( .A1(n767), .A2(n765), .ZN(n728) );
  INV_X1 U560 ( .A(n728), .ZN(n733) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n692) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NOR2_X1 U563 ( .A1(G651), .A2(n637), .ZN(n649) );
  INV_X1 U564 ( .A(G2105), .ZN(n516) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n516), .ZN(n567) );
  NAND2_X1 U566 ( .A1(G126), .A2(n567), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT88), .ZN(n520) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n518), .Z(n902) );
  NAND2_X1 U569 ( .A1(n902), .A2(G138), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U571 ( .A1(n516), .A2(G2104), .ZN(n901) );
  NAND2_X1 U572 ( .A1(G102), .A2(n901), .ZN(n523) );
  INV_X1 U573 ( .A(G2104), .ZN(n521) );
  NOR2_X1 U574 ( .A1(n516), .A2(n521), .ZN(n896) );
  NAND2_X1 U575 ( .A1(G114), .A2(n896), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U577 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U578 ( .A(G651), .ZN(n529) );
  NOR2_X1 U579 ( .A1(G543), .A2(n529), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n526), .Z(n647) );
  NAND2_X1 U581 ( .A1(G64), .A2(n647), .ZN(n528) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  NAND2_X1 U583 ( .A1(G52), .A2(n649), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U586 ( .A1(G90), .A2(n653), .ZN(n532) );
  OR2_X1 U587 ( .A1(n529), .A2(n637), .ZN(n530) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(n530), .ZN(n654) );
  NAND2_X1 U589 ( .A1(G77), .A2(n654), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U591 ( .A(KEYINPUT70), .B(n533), .Z(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT9), .B(n534), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(G171) );
  XOR2_X1 U594 ( .A(G2435), .B(G2427), .Z(n538) );
  XNOR2_X1 U595 ( .A(G2446), .B(G2454), .ZN(n537) );
  XNOR2_X1 U596 ( .A(n538), .B(n537), .ZN(n544) );
  XOR2_X1 U597 ( .A(G2451), .B(G2430), .Z(n540) );
  XNOR2_X1 U598 ( .A(G1348), .B(G1341), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U600 ( .A(G2438), .B(G2443), .Z(n541) );
  XNOR2_X1 U601 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U602 ( .A(n544), .B(n543), .Z(n545) );
  AND2_X1 U603 ( .A1(G14), .A2(n545), .ZN(G401) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U605 ( .A1(G111), .A2(n896), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G135), .A2(n902), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n551) );
  INV_X1 U608 ( .A(n567), .ZN(n548) );
  INV_X1 U609 ( .A(n548), .ZN(n897) );
  NAND2_X1 U610 ( .A1(n897), .A2(G123), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT18), .B(n549), .Z(n550) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n901), .A2(G99), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n1003) );
  XNOR2_X1 U615 ( .A(G2096), .B(n1003), .ZN(n554) );
  OR2_X1 U616 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U617 ( .A(G69), .ZN(G235) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(G88), .A2(n653), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G75), .A2(n654), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G62), .A2(n647), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G50), .A2(n649), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(G166) );
  INV_X1 U627 ( .A(KEYINPUT23), .ZN(n563) );
  AND2_X1 U628 ( .A1(n516), .A2(G101), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G2104), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT66), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G137), .A2(n902), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G113), .A2(n896), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G125), .A2(n567), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(G160) );
  NAND2_X1 U638 ( .A1(G89), .A2(n653), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT77), .B(n572), .Z(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G76), .A2(n654), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT5), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G63), .A2(n647), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G51), .A2(n649), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U653 ( .A(G223), .ZN(n843) );
  NAND2_X1 U654 ( .A1(n843), .A2(G567), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U656 ( .A1(G81), .A2(n653), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n585), .B(KEYINPUT12), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT72), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G68), .A2(n654), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(n589), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G56), .A2(n647), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n590), .Z(n593) );
  NAND2_X1 U664 ( .A1(G43), .A2(n649), .ZN(n591) );
  XNOR2_X1 U665 ( .A(KEYINPUT73), .B(n591), .ZN(n592) );
  NOR2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n929) );
  INV_X1 U668 ( .A(G860), .ZN(n617) );
  OR2_X1 U669 ( .A1(n929), .A2(n617), .ZN(G153) );
  XOR2_X1 U670 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G54), .A2(n649), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G79), .A2(n654), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n647), .A2(G66), .ZN(n598) );
  XOR2_X1 U676 ( .A(KEYINPUT75), .B(n598), .Z(n600) );
  NAND2_X1 U677 ( .A1(n653), .A2(G92), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n601), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT15), .ZN(n925) );
  INV_X1 U682 ( .A(G868), .ZN(n670) );
  NAND2_X1 U683 ( .A1(n925), .A2(n670), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G91), .A2(n653), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G78), .A2(n654), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT71), .B(n609), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G65), .A2(n647), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G53), .A2(n649), .ZN(n610) );
  AND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G299) );
  NOR2_X1 U693 ( .A1(G868), .A2(G299), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT78), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n670), .A2(G286), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U697 ( .A1(n617), .A2(G559), .ZN(n618) );
  INV_X1 U698 ( .A(n925), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n618), .A2(n624), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U701 ( .A1(G868), .A2(n929), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G868), .A2(n624), .ZN(n620) );
  NOR2_X1 U703 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(n623), .Z(G282) );
  NAND2_X1 U706 ( .A1(n624), .A2(G559), .ZN(n667) );
  XNOR2_X1 U707 ( .A(n929), .B(n667), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n625), .A2(G860), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G93), .A2(n653), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G80), .A2(n654), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G67), .A2(n647), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G55), .A2(n649), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n669) );
  XOR2_X1 U716 ( .A(n632), .B(n669), .Z(G145) );
  NAND2_X1 U717 ( .A1(G49), .A2(n649), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U720 ( .A1(n647), .A2(n635), .ZN(n636) );
  XNOR2_X1 U721 ( .A(n636), .B(KEYINPUT80), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G48), .A2(n649), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G86), .A2(n653), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n654), .A2(G73), .ZN(n642) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(G61), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U732 ( .A1(n647), .A2(G60), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n648), .B(KEYINPUT68), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G47), .A2(n649), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U736 ( .A(KEYINPUT69), .B(n652), .ZN(n658) );
  NAND2_X1 U737 ( .A1(G85), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(G72), .A2(n654), .ZN(n655) );
  AND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G290) );
  INV_X1 U741 ( .A(G299), .ZN(n720) );
  XNOR2_X1 U742 ( .A(n720), .B(n929), .ZN(n662) );
  XNOR2_X1 U743 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U744 ( .A(G305), .B(KEYINPUT82), .ZN(n659) );
  XNOR2_X1 U745 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n662), .B(n661), .ZN(n664) );
  XNOR2_X1 U747 ( .A(G290), .B(G166), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n669), .B(n665), .ZN(n666) );
  XNOR2_X1 U750 ( .A(G288), .B(n666), .ZN(n850) );
  XNOR2_X1 U751 ( .A(n667), .B(n850), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n674), .ZN(n676) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n675) );
  XNOR2_X1 U759 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G2072), .A2(n677), .ZN(G158) );
  XNOR2_X1 U761 ( .A(KEYINPUT84), .B(G44), .ZN(n678) );
  XNOR2_X1 U762 ( .A(n678), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n679) );
  XNOR2_X1 U764 ( .A(KEYINPUT22), .B(n679), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n680), .A2(G96), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n681), .A2(G218), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n682), .B(KEYINPUT85), .ZN(n848) );
  NAND2_X1 U768 ( .A1(n848), .A2(G2106), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G120), .A2(G108), .ZN(n683) );
  NOR2_X1 U770 ( .A1(G235), .A2(n683), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n684), .A2(G57), .ZN(n685) );
  XNOR2_X1 U772 ( .A(n685), .B(KEYINPUT86), .ZN(n849) );
  NAND2_X1 U773 ( .A1(G567), .A2(n849), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n924) );
  NAND2_X1 U775 ( .A1(G661), .A2(G483), .ZN(n688) );
  XOR2_X1 U776 ( .A(KEYINPUT87), .B(n688), .Z(n689) );
  NOR2_X1 U777 ( .A1(n924), .A2(n689), .ZN(n846) );
  NAND2_X1 U778 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  NOR2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n797) );
  NOR2_X1 U781 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U782 ( .A1(n797), .A2(n690), .ZN(n942) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n767) );
  INV_X1 U784 ( .A(KEYINPUT64), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n692), .B(n691), .ZN(n765) );
  INV_X1 U786 ( .A(G1996), .ZN(n976) );
  NOR2_X1 U787 ( .A1(n733), .A2(n976), .ZN(n694) );
  XOR2_X1 U788 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n693) );
  XNOR2_X1 U789 ( .A(n694), .B(n693), .ZN(n697) );
  AND2_X1 U790 ( .A1(n733), .A2(G1341), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n695), .A2(n929), .ZN(n696) );
  XNOR2_X1 U792 ( .A(n698), .B(KEYINPUT65), .ZN(n709) );
  NOR2_X1 U793 ( .A1(n925), .A2(n709), .ZN(n699) );
  XNOR2_X1 U794 ( .A(n699), .B(KEYINPUT97), .ZN(n708) );
  NAND2_X1 U795 ( .A1(G2067), .A2(n728), .ZN(n702) );
  NAND2_X1 U796 ( .A1(KEYINPUT98), .A2(KEYINPUT99), .ZN(n700) );
  NOR2_X1 U797 ( .A1(n702), .A2(n700), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n733), .A2(G1348), .ZN(n701) );
  XNOR2_X1 U799 ( .A(KEYINPUT98), .B(n701), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U801 ( .A1(KEYINPUT99), .A2(n704), .ZN(n705) );
  NOR2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n717) );
  NAND2_X1 U804 ( .A1(n925), .A2(n709), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n728), .A2(G2072), .ZN(n710) );
  XNOR2_X1 U806 ( .A(n710), .B(KEYINPUT27), .ZN(n712) );
  INV_X1 U807 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U808 ( .A1(n949), .A2(n728), .ZN(n711) );
  NOR2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n719) );
  NOR2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n714) );
  XNOR2_X1 U811 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n713) );
  XNOR2_X1 U812 ( .A(n714), .B(n713), .ZN(n718) );
  AND2_X1 U813 ( .A1(n715), .A2(n718), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n724) );
  INV_X1 U815 ( .A(n718), .ZN(n722) );
  NAND2_X1 U816 ( .A1(n720), .A2(n719), .ZN(n721) );
  OR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n726) );
  OR2_X1 U819 ( .A1(n728), .A2(G1961), .ZN(n730) );
  XNOR2_X1 U820 ( .A(G2078), .B(KEYINPUT25), .ZN(n727) );
  XNOR2_X1 U821 ( .A(n727), .B(KEYINPUT94), .ZN(n979) );
  NAND2_X1 U822 ( .A1(n728), .A2(n979), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n738), .A2(G171), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U826 ( .A1(G8), .A2(n733), .ZN(n815) );
  NOR2_X1 U827 ( .A1(G1966), .A2(n815), .ZN(n757) );
  NOR2_X1 U828 ( .A1(n733), .A2(G2084), .ZN(n758) );
  XNOR2_X1 U829 ( .A(n758), .B(KEYINPUT93), .ZN(n734) );
  NAND2_X1 U830 ( .A1(G8), .A2(n734), .ZN(n735) );
  NOR2_X1 U831 ( .A1(n757), .A2(n735), .ZN(n736) );
  XOR2_X1 U832 ( .A(KEYINPUT30), .B(n736), .Z(n737) );
  NOR2_X1 U833 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U834 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U836 ( .A(KEYINPUT31), .B(n741), .Z(n742) );
  NAND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U838 ( .A1(G286), .A2(G8), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n755), .A2(n745), .ZN(n752) );
  INV_X1 U840 ( .A(G8), .ZN(n750) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n733), .ZN(n747) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n815), .ZN(n746) );
  NOR2_X1 U843 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U844 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U847 ( .A(KEYINPUT101), .B(n755), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT93), .B(n758), .Z(n759) );
  NAND2_X1 U850 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n807) );
  NAND2_X1 U853 ( .A1(n942), .A2(n807), .ZN(n764) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n938) );
  NAND2_X1 U855 ( .A1(n764), .A2(n938), .ZN(n802) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n926) );
  INV_X1 U857 ( .A(n765), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n838) );
  XNOR2_X1 U859 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U860 ( .A1(n838), .A2(n944), .ZN(n818) );
  AND2_X1 U861 ( .A1(n926), .A2(n818), .ZN(n796) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n836) );
  NAND2_X1 U863 ( .A1(G104), .A2(n901), .ZN(n769) );
  NAND2_X1 U864 ( .A1(G140), .A2(n902), .ZN(n768) );
  NAND2_X1 U865 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U866 ( .A(KEYINPUT34), .B(n770), .ZN(n776) );
  NAND2_X1 U867 ( .A1(G116), .A2(n896), .ZN(n772) );
  NAND2_X1 U868 ( .A1(G128), .A2(n897), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U870 ( .A(KEYINPUT89), .B(n773), .ZN(n774) );
  XNOR2_X1 U871 ( .A(KEYINPUT35), .B(n774), .ZN(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n777), .ZN(n914) );
  NOR2_X1 U874 ( .A1(n836), .A2(n914), .ZN(n778) );
  XNOR2_X1 U875 ( .A(n778), .B(KEYINPUT90), .ZN(n1017) );
  NAND2_X1 U876 ( .A1(n838), .A2(n1017), .ZN(n834) );
  NAND2_X1 U877 ( .A1(G105), .A2(n901), .ZN(n779) );
  XNOR2_X1 U878 ( .A(n779), .B(KEYINPUT38), .ZN(n786) );
  NAND2_X1 U879 ( .A1(G141), .A2(n902), .ZN(n781) );
  NAND2_X1 U880 ( .A1(G129), .A2(n897), .ZN(n780) );
  NAND2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n896), .A2(G117), .ZN(n782) );
  XOR2_X1 U883 ( .A(KEYINPUT92), .B(n782), .Z(n783) );
  NOR2_X1 U884 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n913) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n913), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G107), .A2(n896), .ZN(n788) );
  NAND2_X1 U888 ( .A1(G131), .A2(n902), .ZN(n787) );
  NAND2_X1 U889 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U890 ( .A1(G95), .A2(n901), .ZN(n789) );
  XNOR2_X1 U891 ( .A(KEYINPUT91), .B(n789), .ZN(n790) );
  NOR2_X1 U892 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U893 ( .A1(n897), .A2(G119), .ZN(n792) );
  NAND2_X1 U894 ( .A1(n793), .A2(n792), .ZN(n882) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n882), .ZN(n794) );
  NAND2_X1 U896 ( .A1(n795), .A2(n794), .ZN(n1006) );
  NAND2_X1 U897 ( .A1(n838), .A2(n1006), .ZN(n830) );
  AND2_X1 U898 ( .A1(n834), .A2(n830), .ZN(n823) );
  NAND2_X1 U899 ( .A1(n796), .A2(n823), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U901 ( .A1(n815), .A2(n798), .ZN(n799) );
  OR2_X1 U902 ( .A1(n800), .A2(n799), .ZN(n803) );
  OR2_X1 U903 ( .A1(n815), .A2(n803), .ZN(n801) );
  NOR2_X1 U904 ( .A1(n802), .A2(n801), .ZN(n806) );
  INV_X1 U905 ( .A(n803), .ZN(n804) );
  AND2_X1 U906 ( .A1(n804), .A2(KEYINPUT33), .ZN(n805) );
  NOR2_X1 U907 ( .A1(n806), .A2(n805), .ZN(n825) );
  INV_X1 U908 ( .A(n807), .ZN(n813) );
  NAND2_X1 U909 ( .A1(G166), .A2(G8), .ZN(n808) );
  NOR2_X1 U910 ( .A1(G2090), .A2(n808), .ZN(n811) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n809) );
  XOR2_X1 U912 ( .A(n809), .B(KEYINPUT24), .Z(n810) );
  NOR2_X1 U913 ( .A1(n815), .A2(n810), .ZN(n814) );
  OR2_X1 U914 ( .A1(n811), .A2(n814), .ZN(n812) );
  NOR2_X1 U915 ( .A1(n813), .A2(n812), .ZN(n821) );
  INV_X1 U916 ( .A(n814), .ZN(n817) );
  INV_X1 U917 ( .A(n815), .ZN(n816) );
  NAND2_X1 U918 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(KEYINPUT103), .ZN(n841) );
  NOR2_X1 U924 ( .A1(n882), .A2(G1991), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n827), .B(KEYINPUT105), .ZN(n1007) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n828) );
  XOR2_X1 U927 ( .A(n828), .B(KEYINPUT104), .Z(n829) );
  NAND2_X1 U928 ( .A1(n1007), .A2(n829), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n831), .A2(n830), .ZN(n832) );
  OR2_X1 U930 ( .A1(n913), .A2(G1996), .ZN(n1009) );
  NAND2_X1 U931 ( .A1(n832), .A2(n1009), .ZN(n833) );
  XOR2_X1 U932 ( .A(KEYINPUT39), .B(n833), .Z(n835) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n914), .A2(n836), .ZN(n1014) );
  NAND2_X1 U935 ( .A1(n837), .A2(n1014), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U941 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT106), .B(n845), .ZN(n847) );
  NAND2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G188) );
  XNOR2_X1 U945 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XNOR2_X1 U946 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  NOR2_X1 U949 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U951 ( .A(n925), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(G286), .B(G171), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  NOR2_X1 U954 ( .A1(G37), .A2(n853), .ZN(G397) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2090), .B(KEYINPUT108), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n856), .B(G2678), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2100), .Z(n860) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U965 ( .A(G1956), .B(G1961), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1986), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U968 ( .A(G1976), .B(G1981), .Z(n866) );
  XNOR2_X1 U969 ( .A(G1971), .B(G1966), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U972 ( .A(G2474), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n872) );
  XOR2_X1 U974 ( .A(G1991), .B(KEYINPUT109), .Z(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G100), .A2(n901), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G112), .A2(n896), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G124), .A2(n897), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n875), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G136), .A2(n902), .ZN(n876) );
  XNOR2_X1 U982 ( .A(n876), .B(KEYINPUT110), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U984 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U985 ( .A(G160), .B(G164), .Z(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n912) );
  NAND2_X1 U987 ( .A1(G118), .A2(n896), .ZN(n884) );
  NAND2_X1 U988 ( .A1(G130), .A2(n897), .ZN(n883) );
  NAND2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U990 ( .A(KEYINPUT111), .B(n885), .Z(n890) );
  NAND2_X1 U991 ( .A1(G106), .A2(n901), .ZN(n887) );
  NAND2_X1 U992 ( .A1(G142), .A2(n902), .ZN(n886) );
  NAND2_X1 U993 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U994 ( .A(n888), .B(KEYINPUT45), .Z(n889) );
  NOR2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n891), .B(n1003), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n893) );
  XNOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n892) );
  XNOR2_X1 U999 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U1000 ( .A(n895), .B(n894), .Z(n910) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n896), .ZN(n899) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U1003 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1004 ( .A(n900), .B(KEYINPUT47), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n901), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n902), .ZN(n903) );
  NAND2_X1 U1007 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1008 ( .A(KEYINPUT114), .B(n905), .Z(n906) );
  NAND2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(n908), .B(KEYINPUT115), .ZN(n999) );
  XNOR2_X1 U1011 ( .A(G162), .B(n999), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1014 ( .A(n914), .B(n913), .Z(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n917), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n924), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(G397), .A2(n919), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n922), .A2(G395), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n923), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1024 ( .A(G308), .ZN(G225) );
  INV_X1 U1025 ( .A(n924), .ZN(G319) );
  INV_X1 U1026 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1027 ( .A(KEYINPUT56), .B(G16), .ZN(n948) );
  XNOR2_X1 U1028 ( .A(G1348), .B(n925), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G168), .B(G1966), .ZN(n927) );
  NAND2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(n928), .B(KEYINPUT57), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G1341), .B(KEYINPUT122), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n930), .B(n929), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1040 ( .A(G171), .B(G1961), .Z(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n1030) );
  XOR2_X1 U1046 ( .A(G1341), .B(G19), .Z(n951) );
  XNOR2_X1 U1047 ( .A(n949), .B(G20), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G1981), .B(G6), .Z(n955) );
  XOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT123), .Z(n952) );
  XNOR2_X1 U1051 ( .A(G4), .B(n952), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(n953), .B(KEYINPUT59), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT60), .B(n958), .Z(n960) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G21), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT124), .B(n961), .Z(n963) );
  XNOR2_X1 U1059 ( .A(G1961), .B(G5), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT125), .B(n964), .ZN(n972) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n970) );
  XOR2_X1 U1063 ( .A(G1986), .B(G24), .Z(n968) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1068 ( .A(n970), .B(n969), .Z(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT61), .B(n973), .Z(n974) );
  NOR2_X1 U1071 ( .A1(G16), .A2(n974), .ZN(n975) );
  XOR2_X1 U1072 ( .A(KEYINPUT127), .B(n975), .Z(n1028) );
  XOR2_X1 U1073 ( .A(KEYINPUT120), .B(G29), .Z(n996) );
  XNOR2_X1 U1074 ( .A(G1991), .B(G25), .ZN(n986) );
  XOR2_X1 U1075 ( .A(G2067), .B(G26), .Z(n978) );
  XNOR2_X1 U1076 ( .A(n976), .B(G32), .ZN(n977) );
  NAND2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n983) );
  XOR2_X1 U1078 ( .A(G2072), .B(G33), .Z(n981) );
  XNOR2_X1 U1079 ( .A(n979), .B(G27), .ZN(n980) );
  NAND2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1082 ( .A(KEYINPUT119), .B(n984), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(G28), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n988), .B(KEYINPUT53), .ZN(n991) );
  XOR2_X1 U1086 ( .A(G2084), .B(G34), .Z(n989) );
  XNOR2_X1 U1087 ( .A(KEYINPUT54), .B(n989), .ZN(n990) );
  NAND2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1089 ( .A(G35), .B(G2090), .ZN(n992) );
  NOR2_X1 U1090 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1091 ( .A(KEYINPUT55), .B(n994), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1093 ( .A1(n997), .A2(G11), .ZN(n998) );
  XNOR2_X1 U1094 ( .A(n998), .B(KEYINPUT121), .ZN(n1026) );
  XOR2_X1 U1095 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1002), .Z(n1020) );
  XNOR2_X1 U1099 ( .A(G160), .B(G2084), .ZN(n1004) );
  NAND2_X1 U1100 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1101 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1102 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G162), .B(G2090), .ZN(n1010) );
  NAND2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1105 ( .A(KEYINPUT51), .B(n1011), .Z(n1012) );
  NOR2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1109 ( .A(KEYINPUT118), .B(n1018), .Z(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  INV_X1 U1112 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

