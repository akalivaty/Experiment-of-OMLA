//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT66), .A2(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT66), .A2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(G119), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n200), .B1(new_n203), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n207), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT23), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT73), .B(G110), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n203), .A2(new_n208), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT24), .B(G110), .Z(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n199), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT74), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n199), .B(new_n220), .C1(new_n214), .C2(new_n217), .ZN(new_n221));
  OAI21_X1  g035(.A(G110), .B1(new_n209), .B2(new_n212), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT71), .B(G110), .C1(new_n209), .C2(new_n212), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n227));
  INV_X1    g041(.A(new_n196), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n196), .A2(KEYINPUT72), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n230), .A2(new_n231), .B1(new_n215), .B2(new_n216), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n219), .A2(new_n221), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT75), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT22), .B(G137), .Z(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n188), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n221), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n226), .A2(new_n232), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT76), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n244), .A3(new_n238), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n239), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n189), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(new_n239), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n250), .ZN(new_n252));
  OAI22_X1  g066(.A1(new_n248), .A2(new_n251), .B1(new_n189), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT32), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n197), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n201), .A2(new_n202), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n264), .A3(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n255), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n268));
  AOI22_X1  g082(.A1(new_n268), .A2(new_n257), .B1(new_n201), .B2(new_n202), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT68), .B(new_n265), .C1(new_n269), .C2(new_n256), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G137), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(G137), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n271), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .A4(new_n272), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n267), .A2(new_n270), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n204), .A2(G116), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT67), .B(G119), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(G116), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT2), .B(G113), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n277), .A2(new_n279), .A3(new_n272), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n256), .A2(KEYINPUT0), .A3(G128), .ZN(new_n297));
  INV_X1    g111(.A(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G146), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n257), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  OR2_X1    g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n296), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n284), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n234), .A3(G210), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT27), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G101), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n284), .A2(KEYINPUT30), .A3(new_n304), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n313));
  INV_X1    g127(.A(new_n263), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n282), .B1(new_n314), .B2(new_n265), .ZN(new_n315));
  INV_X1    g129(.A(new_n304), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n317), .A3(new_n292), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n311), .A2(KEYINPUT31), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT31), .B1(new_n311), .B2(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n305), .A2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n284), .A2(new_n322), .A3(new_n293), .A4(new_n304), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n315), .A2(new_n316), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n321), .A2(new_n323), .B1(new_n292), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n310), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n319), .A2(new_n320), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT70), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n254), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n254), .A3(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n321), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(new_n292), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n327), .A2(KEYINPUT29), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n284), .A2(new_n304), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n321), .A2(new_n323), .B1(new_n292), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n310), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n318), .A2(new_n305), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n343), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G472), .B1(new_n347), .B2(G902), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n253), .B1(new_n336), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT101), .ZN(new_n351));
  XNOR2_X1  g165(.A(G113), .B(G122), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(G104), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n353), .B(KEYINPUT93), .Z(new_n354));
  NAND2_X1  g168(.A1(new_n191), .A2(new_n193), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT92), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(G146), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n198), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n306), .A2(new_n234), .A3(G214), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n298), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n306), .A2(new_n234), .A3(G143), .A4(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT18), .A2(G131), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(new_n364), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI211_X1 g183(.A(KEYINPUT91), .B(new_n364), .C1(new_n362), .C2(new_n363), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n360), .B(new_n365), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(G131), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n280), .A3(new_n363), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT94), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n372), .A2(KEYINPUT94), .A3(new_n373), .A4(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n367), .A2(KEYINPUT17), .A3(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n230), .A2(new_n231), .A3(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n354), .B(new_n371), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n357), .A2(KEYINPUT19), .A3(new_n358), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n355), .A2(KEYINPUT19), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n197), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n374), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n196), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n371), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n353), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT20), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n394), .A3(new_n391), .ZN(new_n395));
  INV_X1    g209(.A(new_n353), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n230), .A2(new_n231), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n397), .A2(new_n380), .A3(new_n377), .A4(new_n378), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n398), .B2(new_n371), .ZN(new_n399));
  INV_X1    g213(.A(new_n382), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n188), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n393), .A2(new_n395), .B1(new_n401), .B2(G475), .ZN(new_n402));
  NAND2_X1  g216(.A1(G234), .A2(G237), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(G952), .A3(new_n234), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(G902), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT21), .B(G898), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT9), .B(G234), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n412), .A2(new_n187), .A3(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT98), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n201), .A2(G143), .A3(new_n202), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n298), .A2(G128), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n271), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n271), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n418), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G134), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT97), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT79), .B(G107), .ZN(new_n427));
  INV_X1    g241(.A(G116), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G122), .ZN(new_n429));
  INV_X1    g243(.A(G122), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT95), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(G116), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(G122), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT95), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n427), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OR3_X1    g251(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT14), .ZN(new_n438));
  INV_X1    g252(.A(G107), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n431), .B2(KEYINPUT14), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n417), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n421), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT13), .A2(G134), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n417), .A2(new_n418), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n435), .B1(new_n433), .B2(new_n434), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT79), .A2(G107), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT79), .A2(G107), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n444), .B(new_n446), .C1(new_n452), .C2(new_n437), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT96), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n432), .A2(new_n427), .A3(new_n436), .ZN(new_n456));
  INV_X1    g270(.A(new_n423), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n455), .A2(new_n456), .B1(new_n457), .B2(new_n445), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT96), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n444), .ZN(new_n460));
  AOI221_X4 g274(.A(new_n415), .B1(new_n426), .B2(new_n441), .C1(new_n454), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n460), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n426), .A2(new_n441), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n414), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT100), .B(new_n188), .C1(new_n461), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n453), .A2(KEYINPUT96), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n459), .B1(new_n458), .B2(new_n444), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n415), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n463), .A3(new_n414), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n470), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n477), .A2(KEYINPUT100), .A3(new_n188), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n351), .B1(new_n411), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n480), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(KEYINPUT101), .A3(new_n402), .A4(new_n410), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  INV_X1    g301(.A(G104), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT3), .ZN(new_n489));
  OR2_X1    g303(.A1(KEYINPUT79), .A2(G107), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT79), .A2(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n439), .B1(new_n493), .B2(G104), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(G104), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n487), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n495), .A2(new_n449), .A3(new_n450), .ZN(new_n501));
  AOI21_X1  g315(.A(G107), .B1(new_n488), .B2(KEYINPUT3), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n489), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(G101), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n496), .A3(new_n487), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n497), .A2(new_n500), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n292), .B(new_n499), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n492), .A2(new_n496), .A3(new_n487), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n488), .B1(new_n449), .B2(new_n450), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n427), .A2(KEYINPUT82), .A3(new_n488), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT81), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(G104), .B2(new_n439), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n488), .A2(KEYINPUT81), .A3(G107), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n509), .B1(new_n518), .B2(G101), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n205), .A2(new_n207), .A3(new_n520), .A4(G116), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n521), .A2(G113), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n428), .A2(G119), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT5), .B(new_n523), .C1(new_n210), .C2(new_n428), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n522), .A2(new_n524), .B1(new_n287), .B2(new_n289), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n519), .A2(KEYINPUT87), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT87), .B1(new_n519), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G110), .B(G122), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n529), .B(new_n508), .C1(new_n526), .C2(new_n527), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n518), .A2(G101), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n535), .A3(new_n505), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n519), .A2(KEYINPUT87), .A3(new_n525), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n540), .B2(new_n508), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n543), .A3(new_n530), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n533), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n192), .B(new_n265), .C1(new_n269), .C2(new_n256), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n303), .A2(new_n297), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G125), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n234), .A2(G224), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G210), .B1(G237), .B2(G902), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n548), .A2(KEYINPUT7), .A3(new_n552), .A4(new_n550), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n548), .A2(new_n550), .B1(KEYINPUT7), .B2(new_n552), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(KEYINPUT90), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(KEYINPUT90), .B2(new_n558), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n529), .B(KEYINPUT8), .Z(new_n561));
  OR2_X1    g375(.A1(new_n519), .A2(new_n525), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n536), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI211_X1 g379(.A(KEYINPUT89), .B(new_n561), .C1(new_n562), .C2(new_n536), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n560), .B(new_n532), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n188), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n555), .A2(new_n556), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n556), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n545), .B(new_n544), .C1(new_n534), .C2(new_n541), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n553), .B1(new_n572), .B2(new_n533), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n573), .B2(new_n568), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n486), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G221), .B1(new_n412), .B2(G902), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT77), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n519), .A2(new_n267), .A3(new_n270), .A4(KEYINPUT10), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n549), .B1(new_n498), .B2(new_n497), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n506), .B2(new_n507), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT84), .ZN(new_n583));
  INV_X1    g397(.A(new_n296), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n300), .A2(new_n211), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n265), .B(new_n585), .C1(new_n258), .C2(new_n299), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n535), .A2(new_n505), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n579), .A3(new_n584), .A4(new_n581), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT84), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n519), .A2(new_n263), .A3(new_n266), .ZN(new_n594));
  INV_X1    g408(.A(new_n587), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n296), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT12), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(KEYINPUT12), .B(new_n296), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n234), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT78), .ZN(new_n602));
  XNOR2_X1  g416(.A(G110), .B(G140), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n589), .A2(new_n581), .A3(new_n579), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n296), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT86), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n610), .A3(new_n296), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n609), .A2(new_n611), .B1(new_n590), .B2(new_n592), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n606), .B1(new_n612), .B2(new_n605), .ZN(new_n613));
  INV_X1    g427(.A(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n188), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n600), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n604), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT85), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n591), .A2(KEYINPUT84), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n591), .A2(KEYINPUT84), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n618), .B(new_n605), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n609), .A2(new_n611), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n604), .B1(new_n590), .B2(new_n592), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n618), .ZN(new_n625));
  OAI211_X1 g439(.A(G469), .B(new_n617), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n614), .A2(new_n188), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n615), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n484), .A2(new_n575), .A3(new_n578), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n350), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n487), .ZN(G3));
  AND2_X1   g446(.A1(new_n629), .A2(new_n578), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n556), .B1(new_n555), .B2(new_n569), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n573), .A2(new_n571), .A3(new_n568), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n485), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n409), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT31), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n312), .A2(new_n317), .A3(new_n292), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n305), .A2(new_n310), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n311), .A2(KEYINPUT31), .A3(new_n318), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n337), .A2(new_n338), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n327), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n644), .B2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n329), .A2(new_n332), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n253), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n461), .B2(new_n464), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n477), .A2(KEYINPUT102), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n475), .A2(KEYINPUT33), .A3(new_n476), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT103), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n475), .A2(new_n657), .A3(KEYINPUT33), .A4(new_n476), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n466), .A2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n654), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n477), .A2(new_n188), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n466), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n402), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AND4_X1   g478(.A1(new_n633), .A2(new_n637), .A3(new_n648), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT104), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND3_X1  g482(.A1(new_n480), .A2(new_n402), .A3(new_n410), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT105), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n633), .A2(new_n575), .A3(new_n648), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n238), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n233), .B(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n189), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n188), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n248), .B2(new_n251), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n681), .B(new_n684), .C1(new_n248), .C2(new_n251), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n646), .A3(new_n645), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n630), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NOR3_X1   g503(.A1(new_n644), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n348), .B1(new_n690), .B2(new_n333), .ZN(new_n691));
  INV_X1    g505(.A(new_n402), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n404), .B(KEYINPUT107), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n694), .B1(new_n695), .B2(new_n407), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n482), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n683), .A2(new_n691), .A3(new_n685), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n575), .A2(new_n578), .A3(new_n629), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n211), .ZN(G30));
  XOR2_X1   g515(.A(new_n696), .B(KEYINPUT39), .Z(new_n702));
  NAND3_X1  g516(.A1(new_n633), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n629), .A2(new_n578), .ZN(new_n705));
  INV_X1    g519(.A(new_n702), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n710), .B1(new_n703), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n570), .A2(new_n574), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n682), .A2(new_n482), .A3(new_n402), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n341), .A2(new_n292), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n328), .B1(new_n716), .B2(new_n305), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n318), .B2(new_n311), .ZN(new_n718));
  OAI21_X1  g532(.A(G472), .B1(new_n718), .B2(G902), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n690), .B2(new_n333), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n714), .A2(new_n485), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  AOI211_X1 g538(.A(new_n402), .B(new_n696), .C1(new_n661), .C2(new_n663), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n683), .A3(new_n691), .A4(new_n685), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n699), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n197), .ZN(G48));
  AOI21_X1  g542(.A(new_n610), .B1(new_n607), .B2(new_n296), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n607), .A2(new_n610), .A3(new_n296), .ZN(new_n730));
  OAI22_X1  g544(.A1(new_n729), .A2(new_n730), .B1(new_n619), .B2(new_n620), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n731), .A2(new_n604), .B1(new_n600), .B2(new_n624), .ZN(new_n732));
  OAI21_X1  g546(.A(G469), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n578), .A3(new_n615), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n637), .A2(new_n349), .A3(new_n664), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND4_X1  g552(.A1(new_n349), .A2(new_n735), .A3(new_n670), .A4(new_n575), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND4_X1  g554(.A1(new_n484), .A2(new_n683), .A3(new_n691), .A4(new_n685), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n636), .B2(new_n734), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n732), .A2(G469), .A3(G902), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n614), .B1(new_n613), .B2(new_n188), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n575), .A3(KEYINPUT109), .A4(new_n578), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n741), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n204), .ZN(G21));
  NOR2_X1   g563(.A1(new_n482), .A2(new_n402), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n575), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n319), .A2(new_n320), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n342), .A2(new_n328), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n332), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n645), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n253), .A2(new_n755), .A3(new_n409), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n751), .A2(new_n735), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  INV_X1    g572(.A(new_n251), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n678), .B1(new_n252), .B2(KEYINPUT25), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n680), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n725), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n743), .B2(new_n747), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n192), .ZN(G27));
  NAND3_X1  g579(.A1(new_n570), .A2(new_n574), .A3(new_n485), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n633), .A2(new_n349), .A3(new_n725), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n705), .A2(new_n766), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT42), .A3(new_n349), .A4(new_n725), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NAND3_X1  g588(.A1(new_n767), .A2(new_n578), .A3(new_n629), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n350), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n697), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  OAI21_X1  g592(.A(new_n617), .B1(new_n623), .B2(new_n625), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n614), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n628), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n744), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n628), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n578), .A3(new_n702), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n791), .A3(new_n578), .A4(new_n702), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n692), .B1(new_n661), .B2(new_n663), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT43), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n795), .A2(new_n647), .A3(new_n682), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n766), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n790), .A2(new_n792), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  INV_X1    g619(.A(new_n696), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n664), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n253), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n807), .A2(new_n766), .A3(new_n691), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n788), .B2(new_n578), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n811), .B(new_n577), .C1(new_n786), .C2(new_n787), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(new_n714), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n746), .B(KEYINPUT49), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n808), .A2(new_n578), .A3(new_n485), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n720), .A3(new_n794), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n699), .B1(new_n726), .B2(new_n698), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n720), .A2(new_n761), .A3(new_n806), .A4(new_n750), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n699), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n764), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n824), .B2(KEYINPUT52), .ZN(new_n825));
  INV_X1    g639(.A(new_n821), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n743), .A2(new_n747), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n807), .A2(new_n761), .A3(new_n755), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n823), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n826), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n770), .A2(new_n772), .B1(new_n776), .B2(new_n697), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n482), .A2(new_n692), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n664), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n637), .A2(new_n633), .A3(new_n648), .A4(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n736), .A2(new_n840), .A3(new_n757), .A4(new_n739), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n630), .B1(new_n350), .B2(new_n686), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n748), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n692), .A2(new_n480), .A3(new_n696), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n683), .A2(new_n691), .A3(new_n685), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n775), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n775), .B2(new_n763), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n828), .A2(new_n771), .A3(KEYINPUT112), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n837), .A2(new_n841), .A3(new_n843), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n836), .B2(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n764), .A2(new_n821), .A3(new_n832), .A4(new_n823), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n834), .B2(new_n826), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n837), .A2(new_n841), .A3(new_n843), .A4(new_n850), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n851), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n795), .A2(new_n798), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n253), .A2(new_n755), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n694), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n766), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n810), .A2(new_n812), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n744), .A2(new_n745), .A3(new_n578), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n867), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n815), .A2(new_n486), .A3(new_n735), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT50), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n877), .B1(new_n881), .B2(KEYINPUT116), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n867), .B2(new_n875), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n734), .A2(new_n766), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n720), .A2(new_n253), .A3(new_n404), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n661), .A2(new_n402), .A3(new_n663), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n865), .A2(new_n694), .A3(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(new_n762), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n883), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n873), .A2(KEYINPUT51), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT51), .B1(new_n873), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n888), .A2(new_n350), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT48), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n885), .A3(new_n664), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G952), .A3(new_n234), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n874), .B2(new_n827), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n864), .A2(new_n892), .A3(new_n893), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(G952), .A2(G953), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT117), .Z(new_n902));
  OAI21_X1  g716(.A(new_n819), .B1(new_n900), .B2(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n547), .B(KEYINPUT118), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n553), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n860), .A2(new_n862), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(G902), .ZN(new_n910));
  INV_X1    g724(.A(G210), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n904), .B(new_n908), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n234), .A2(G952), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT119), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n907), .ZN(G51));
  INV_X1    g731(.A(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n863), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n627), .B(KEYINPUT57), .Z(new_n921));
  OAI21_X1  g735(.A(new_n613), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n188), .B1(new_n860), .B2(new_n862), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(new_n781), .A3(new_n782), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n918), .B1(new_n922), .B2(new_n924), .ZN(G54));
  AND3_X1   g739(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n390), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(G60));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n466), .A2(new_n188), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n835), .B1(new_n854), .B2(KEYINPUT113), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n824), .A2(new_n820), .A3(KEYINPUT52), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n851), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n857), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n851), .B(KEYINPUT53), .C1(new_n854), .C2(new_n853), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n861), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n654), .A2(new_n659), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT120), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(KEYINPUT122), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n933), .B1(new_n859), .B2(new_n863), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n919), .A2(new_n863), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n945), .A2(new_n933), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n918), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n946), .A2(new_n949), .A3(new_n952), .ZN(G63));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT60), .Z(new_n956));
  AND2_X1   g770(.A1(new_n909), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n249), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n233), .A2(new_n238), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n914), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n909), .A2(new_n956), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n677), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n954), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n958), .B2(new_n959), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT61), .A4(new_n914), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(G66));
  INV_X1    g782(.A(new_n408), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n234), .B1(new_n969), .B2(G224), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n841), .A2(new_n843), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n234), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n905), .B1(G898), .B2(new_n234), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n839), .A2(new_n349), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n709), .A2(new_n767), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n981), .A2(new_n712), .A3(new_n721), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n764), .A2(new_n821), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n723), .A2(KEYINPUT62), .A3(new_n983), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n804), .A2(new_n813), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n312), .A2(new_n317), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n383), .A2(new_n384), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n976), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n982), .A2(new_n980), .A3(new_n984), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT62), .B1(new_n723), .B2(new_n983), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n978), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n804), .A2(new_n813), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n234), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(KEYINPUT124), .A3(new_n992), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n790), .A2(new_n349), .A3(new_n751), .A4(new_n792), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n837), .A2(new_n983), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n988), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n994), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1007), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n994), .A2(new_n1000), .A3(new_n1009), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G72));
  INV_X1    g825(.A(new_n310), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n345), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n997), .A2(new_n971), .A3(new_n998), .ZN(new_n1014));
  XOR2_X1   g828(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1013), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n345), .A2(new_n1012), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1021), .B(new_n1022), .C1(new_n852), .C2(new_n858), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n971), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n988), .A2(new_n1025), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1026), .A2(new_n1018), .ZN(new_n1027));
  OAI211_X1 g841(.A(KEYINPUT127), .B(new_n914), .C1(new_n1027), .C2(new_n1021), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1021), .B1(new_n1026), .B2(new_n1018), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n918), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1024), .B1(new_n1028), .B2(new_n1031), .ZN(G57));
endmodule


