//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(KEYINPUT74), .A3(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT27), .B(G183gat), .Z(new_n219));
  INV_X1    g018(.A(KEYINPUT28), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G190gat), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT67), .B(G190gat), .Z(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G183gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n223), .B(new_n226), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n222), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT69), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  NOR2_X1   g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n245));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n239), .A2(new_n240), .A3(new_n250), .A4(new_n241), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT24), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n238), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n255), .B(new_n256), .C1(new_n221), .C2(G183gat), .ZN(new_n257));
  AND4_X1   g056(.A1(KEYINPUT25), .A2(new_n245), .A3(new_n246), .A4(new_n248), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n252), .A2(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n237), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(KEYINPUT29), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n231), .A2(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n223), .A2(new_n226), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(new_n267), .B2(new_n222), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n257), .A2(new_n258), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n263), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n218), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT75), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n237), .A2(new_n259), .B1(KEYINPUT29), .B2(new_n261), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n271), .A3(new_n260), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n213), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n218), .ZN(new_n280));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT76), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n274), .A2(new_n277), .A3(new_n280), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n202), .B1(new_n287), .B2(KEYINPUT30), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(KEYINPUT79), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n284), .B(KEYINPUT77), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n288), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OR3_X1    g093(.A1(new_n286), .A2(KEYINPUT78), .A3(new_n289), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT78), .B1(new_n286), .B2(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G141gat), .B(G148gat), .Z(new_n299));
  XNOR2_X1  g098(.A(G155gat), .B(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n306));
  INV_X1    g105(.A(new_n301), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n309), .A2(KEYINPUT80), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(KEYINPUT80), .ZN(new_n311));
  OAI211_X1 g110(.A(KEYINPUT81), .B(new_n301), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n312), .A3(new_n299), .ZN(new_n313));
  INV_X1    g112(.A(new_n300), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n317));
  OAI21_X1  g116(.A(G127gat), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319));
  OAI221_X1 g118(.A(new_n318), .B1(G127gat), .B2(G134gat), .C1(KEYINPUT1), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(KEYINPUT71), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n322), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT1), .ZN(new_n324));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT83), .ZN(new_n330));
  INV_X1    g129(.A(new_n328), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n334), .A3(KEYINPUT4), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT82), .A4(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT82), .B1(new_n328), .B2(KEYINPUT4), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n328), .B2(KEYINPUT4), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT83), .B(new_n332), .C1(new_n315), .C2(new_n327), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n320), .A2(new_n326), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n315), .B2(new_n341), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n336), .B(new_n340), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT39), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n315), .A2(new_n327), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n352), .B2(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(new_n350), .A3(new_n348), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT40), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n347), .C1(new_n343), .C2(new_n345), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n336), .A2(new_n365), .A3(new_n340), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n348), .B1(new_n331), .B2(new_n351), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n328), .B(new_n332), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n347), .B1(new_n343), .B2(new_n345), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT5), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n358), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n360), .B2(new_n361), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n298), .A2(new_n362), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n370), .ZN(new_n375));
  INV_X1    g174(.A(new_n358), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n371), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n275), .A2(new_n276), .A3(new_n218), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT37), .ZN(new_n383));
  INV_X1    g182(.A(new_n213), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n275), .B2(new_n276), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT88), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT37), .A4(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n274), .A2(new_n277), .A3(new_n280), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n292), .A2(KEYINPUT38), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT89), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n390), .A2(new_n396), .A3(new_n392), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n366), .A2(new_n370), .A3(new_n358), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n378), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n291), .A2(KEYINPUT37), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n284), .A3(new_n392), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n287), .B1(new_n402), .B2(KEYINPUT38), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n381), .A2(new_n398), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n217), .B1(new_n342), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT3), .B1(new_n213), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(new_n315), .ZN(new_n411));
  OAI211_X1 g210(.A(G228gat), .B(G233gat), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n413));
  INV_X1    g212(.A(new_n411), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n315), .B2(new_n341), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n414), .B(new_n415), .C1(new_n213), .C2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n413), .B1(new_n412), .B2(new_n417), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n342), .A2(new_n408), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n218), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n415), .B1(new_n410), .B2(new_n315), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n423), .B2(new_n384), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT86), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n407), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n418), .B2(new_n419), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n422), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n406), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n373), .A2(new_n404), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n431), .A2(KEYINPUT87), .A3(new_n434), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT87), .B1(new_n431), .B2(new_n434), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n399), .A2(new_n441), .A3(new_n378), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n399), .B2(new_n378), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n442), .A2(new_n443), .A3(new_n371), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n379), .A2(new_n380), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n294), .B(new_n297), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n327), .B1(new_n237), .B2(new_n259), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n268), .A2(new_n271), .A3(new_n344), .ZN(new_n448));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT72), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n447), .A2(new_n448), .A3(new_n453), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n450), .B1(new_n447), .B2(new_n448), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n449), .B2(KEYINPUT73), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n458), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G15gat), .B(G43gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n458), .B(new_n460), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT33), .B1(new_n452), .B2(new_n454), .ZN(new_n468));
  INV_X1    g267(.A(new_n465), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n466), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n466), .B2(new_n470), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT36), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n440), .A2(new_n446), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n436), .A2(new_n475), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT35), .B1(new_n446), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n473), .B2(new_n474), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n471), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n470), .A3(new_n472), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(KEYINPUT90), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n431), .A2(new_n489), .A3(new_n434), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n381), .B2(new_n400), .ZN(new_n491));
  INV_X1    g290(.A(new_n298), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n437), .A2(new_n479), .B1(new_n481), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT91), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT14), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n499), .B(new_n503), .C1(G29gat), .C2(G36gat), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n506), .A2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n507), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n505), .B(new_n509), .C1(KEYINPUT92), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n501), .A2(KEYINPUT92), .A3(new_n502), .A4(new_n504), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n501), .A2(new_n502), .A3(new_n509), .A4(new_n504), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n514), .C1(new_n507), .C2(new_n510), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n495), .B1(new_n516), .B2(KEYINPUT17), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(KEYINPUT93), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G1gat), .B2(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G8gat), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n524), .B(new_n527), .C1(G1gat), .C2(new_n521), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT94), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n518), .B1(new_n512), .B2(new_n515), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n516), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n529), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n520), .A2(new_n535), .B1(new_n538), .B2(new_n529), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n537), .ZN(new_n544));
  INV_X1    g343(.A(new_n529), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n516), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n537), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n555), .A3(new_n544), .A4(new_n549), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G64gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(G57gat), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT97), .B(new_n563), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(KEYINPUT96), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(G57gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n572), .A2(new_n573), .B1(new_n562), .B2(new_n561), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n574), .B2(KEYINPUT97), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n571), .B(new_n563), .C1(new_n565), .C2(new_n567), .ZN(new_n576));
  INV_X1    g375(.A(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n570), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n529), .B1(KEYINPUT21), .B2(new_n579), .ZN(new_n584));
  OR3_X1    g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n580), .B(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n584), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT20), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT98), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n585), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n585), .B2(new_n587), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT41), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n599), .B(new_n602), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT7), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n610), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n534), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n520), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT100), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n621), .A2(KEYINPUT100), .B1(new_n601), .B2(new_n600), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n538), .B2(new_n617), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n619), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n604), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(new_n622), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n603), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n598), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G120gat), .B(G148gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT104), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT101), .B1(new_n579), .B2(new_n617), .ZN(new_n641));
  INV_X1    g440(.A(new_n616), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n568), .A2(KEYINPUT96), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n577), .A3(new_n576), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n644), .A2(new_n645), .A3(new_n570), .A4(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n579), .A2(new_n617), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n579), .A2(new_n617), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n640), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n638), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n649), .B2(new_n654), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n579), .B2(new_n617), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n639), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n655), .A2(KEYINPUT103), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(KEYINPUT105), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n660), .A2(new_n667), .A3(new_n639), .A4(new_n662), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n656), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n638), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR4_X1   g470(.A1(new_n494), .A2(new_n560), .A3(new_n634), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n444), .A2(new_n445), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  INV_X1    g476(.A(new_n672), .ZN(new_n678));
  OAI21_X1  g477(.A(G8gat), .B1(new_n678), .B2(new_n492), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n672), .A2(new_n298), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n677), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n684), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT106), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(G1325gat));
  NAND2_X1  g487(.A1(new_n476), .A2(new_n478), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n678), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n488), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n678), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n672), .A2(new_n440), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n494), .A2(new_n560), .ZN(new_n697));
  INV_X1    g496(.A(new_n671), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n597), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n633), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n673), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(G29gat), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n627), .A2(new_n632), .A3(KEYINPUT108), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n627), .B2(new_n632), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT109), .B1(new_n494), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n494), .B2(new_n633), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n479), .A2(new_n437), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n481), .A2(new_n493), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n709), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n711), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n699), .A2(new_n560), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n702), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n701), .A2(G36gat), .A3(new_n492), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n492), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(new_n689), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n718), .A2(new_n727), .A3(new_n719), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n691), .A2(G43gat), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n559), .A3(new_n700), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT111), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT110), .B(KEYINPUT47), .C1(new_n729), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(G43gat), .B2(new_n728), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n733), .A2(new_n737), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n440), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n701), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n701), .A2(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n440), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n720), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n743), .B2(new_n744), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n720), .B2(new_n436), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n698), .A2(new_n634), .A3(new_n559), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n715), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(KEYINPUT114), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(KEYINPUT114), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n702), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n566), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n492), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT49), .B(G64gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n764), .B2(new_n767), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n689), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT115), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n759), .A2(new_n773), .A3(new_n760), .A4(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n761), .B2(new_n691), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1334gat));
  NOR2_X1   g581(.A1(new_n761), .A2(new_n746), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g583(.A1(new_n698), .A2(new_n559), .A3(new_n598), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n718), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT117), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n718), .A2(new_n788), .A3(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n673), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT118), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n787), .A2(new_n792), .A3(new_n673), .A4(new_n789), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(G85gat), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n633), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n559), .A2(new_n598), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n715), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT51), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n715), .A2(new_n799), .A3(new_n795), .A4(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n671), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n605), .A3(new_n673), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n794), .A2(new_n803), .ZN(G1336gat));
  NOR3_X1   g603(.A1(new_n801), .A2(G92gat), .A3(new_n492), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(G92gat), .B1(new_n786), .B2(new_n492), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n298), .A3(new_n789), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n809), .B2(G92gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  AOI21_X1  g611(.A(G99gat), .B1(new_n802), .B2(new_n488), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n787), .A2(new_n789), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n727), .A2(G99gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G1338gat));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n440), .A3(new_n789), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n436), .A2(G106gat), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(G106gat), .B1(new_n802), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n798), .A2(new_n671), .A3(new_n800), .A4(new_n818), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n786), .B2(new_n436), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT119), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n819), .A2(new_n820), .B1(new_n824), .B2(new_n825), .ZN(G1339gat));
  NOR2_X1   g625(.A1(new_n706), .A2(new_n707), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n666), .A2(new_n828), .A3(new_n668), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n660), .A2(new_n662), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n640), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n663), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n638), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT55), .A4(new_n638), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n559), .A3(new_n665), .A4(new_n836), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n543), .A2(new_n537), .B1(new_n546), .B2(new_n548), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n554), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n558), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n671), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n827), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n835), .A2(new_n665), .A3(new_n840), .A4(new_n836), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n708), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n597), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n634), .A2(new_n671), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n560), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n560), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n702), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n492), .A2(new_n852), .A3(new_n436), .A4(new_n475), .ZN(new_n853));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n559), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n845), .A2(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n746), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n691), .B1(new_n856), .B2(KEYINPUT121), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n858), .A3(new_n746), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n702), .A2(new_n298), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n560), .A2(new_n322), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n854), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(G120gat), .B1(new_n853), .B2(new_n671), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n671), .A2(G120gat), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n863), .B2(new_n867), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n869), .A3(new_n598), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n860), .A2(new_n597), .A3(new_n862), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(G1342gat));
  NOR3_X1   g671(.A1(new_n633), .A2(new_n317), .A3(new_n316), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT56), .Z(new_n875));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n633), .A3(new_n862), .ZN(new_n876));
  INV_X1    g675(.A(G134gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n727), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n855), .B2(new_n435), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(KEYINPUT123), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n795), .B1(new_n837), .B2(new_n841), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n844), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n851), .B1(new_n884), .B2(new_n598), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(KEYINPUT57), .A3(new_n440), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n881), .B2(KEYINPUT123), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G141gat), .B1(new_n888), .B2(new_n560), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n727), .A2(new_n298), .A3(new_n436), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n852), .A2(new_n890), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n891), .A2(G141gat), .A3(new_n560), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT124), .B(KEYINPUT58), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n889), .A2(new_n896), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1344gat));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n891), .A2(G148gat), .A3(new_n698), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n879), .B(new_n671), .C1(new_n882), .C2(new_n887), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n855), .A2(new_n435), .A3(new_n880), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n843), .A2(new_n633), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n597), .B1(new_n883), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n847), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n440), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n879), .A2(new_n671), .ZN(new_n912));
  OAI21_X1  g711(.A(G148gat), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n899), .B(new_n901), .C1(new_n905), .C2(new_n914), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n902), .A2(new_n904), .B1(new_n913), .B2(KEYINPUT59), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT125), .B1(new_n916), .B2(new_n900), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n888), .B2(new_n597), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n891), .A2(G155gat), .A3(new_n597), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n888), .B2(new_n708), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n891), .A2(G162gat), .A3(new_n633), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n856), .A2(KEYINPUT121), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n492), .A2(new_n673), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n488), .A3(new_n859), .A4(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n857), .A2(KEYINPUT126), .A3(new_n859), .A4(new_n926), .ZN(new_n930));
  AND4_X1   g729(.A1(G169gat), .A2(new_n929), .A3(new_n559), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n673), .B1(new_n845), .B2(new_n851), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n492), .A2(new_n480), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n559), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n931), .A2(new_n936), .ZN(G1348gat));
  NAND3_X1  g736(.A1(new_n929), .A2(new_n671), .A3(new_n930), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G176gat), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n698), .A2(G176gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n934), .B2(new_n940), .ZN(G1349gat));
  NAND3_X1  g740(.A1(new_n929), .A2(new_n598), .A3(new_n930), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G183gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n935), .A2(new_n227), .A3(new_n598), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n935), .A2(new_n223), .A3(new_n827), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n795), .A3(new_n930), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(G190gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n951), .B2(G190gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  NAND3_X1  g754(.A1(new_n689), .A2(new_n298), .A3(new_n435), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT127), .Z(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n932), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n559), .ZN(new_n959));
  INV_X1    g758(.A(new_n911), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n926), .A2(new_n689), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n559), .A2(G197gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  INV_X1    g763(.A(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n958), .A2(new_n965), .A3(new_n671), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  INV_X1    g766(.A(new_n962), .ZN(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n968), .B2(new_n698), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n958), .A2(new_n205), .A3(new_n598), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n962), .A2(new_n598), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  OAI21_X1  g774(.A(G218gat), .B1(new_n968), .B2(new_n633), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n206), .A3(new_n827), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1355gat));
endmodule


