//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n206), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G116), .A2(G270), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n229), .B1(new_n217), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(G68), .B2(G238), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(G77), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n228), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n212), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n215), .B(new_n221), .C1(new_n237), .C2(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n219), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT70), .B(G107), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT75), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT75), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n269), .B2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n258), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G77), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT6), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(new_n225), .A3(G107), .ZN(new_n275));
  XNOR2_X1  g0075(.A(G97), .B(G107), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(new_n210), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n256), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G97), .ZN(new_n283));
  INV_X1    g0083(.A(new_n256), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n282), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n209), .B2(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(G97), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n219), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT4), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n262), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n264), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(new_n233), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT4), .A2(G244), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n264), .A2(new_n294), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G283), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n264), .A2(new_n294), .A3(G250), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n302), .B2(KEYINPUT4), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n292), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT67), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n290), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n289), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n219), .B1(new_n306), .B2(new_n290), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n308), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G41), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n209), .A2(G45), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT5), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(G41), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(G257), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G274), .B1(new_n319), .B2(G41), .ZN(new_n322));
  INV_X1    g0122(.A(new_n317), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT80), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n324), .C1(KEYINPUT5), .C2(new_n315), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT80), .B1(new_n316), .B2(new_n317), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n314), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n304), .A2(new_n305), .A3(new_n321), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n288), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n302), .A2(KEYINPUT4), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G1698), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n299), .A2(new_n300), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n296), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n292), .B1(new_n314), .B2(new_n327), .ZN(new_n335));
  AOI21_X1  g0135(.A(G169), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT81), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n304), .A2(new_n321), .A3(new_n328), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT81), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n288), .A4(new_n329), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(G200), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(G190), .A3(new_n321), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n279), .A4(new_n287), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n337), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT82), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n337), .A2(new_n345), .A3(KEYINPUT82), .A4(new_n342), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n312), .B1(new_n311), .B2(new_n308), .ZN(new_n350));
  AND4_X1   g0150(.A1(new_n312), .A2(new_n307), .A3(new_n289), .A4(new_n308), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n317), .A2(new_n224), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G274), .B2(new_n317), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n233), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n269), .B(new_n356), .C1(G238), .C2(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G116), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n291), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n355), .A2(new_n305), .A3(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n355), .A2(new_n359), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(G169), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT83), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n223), .A2(new_n225), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n257), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n257), .B2(new_n364), .ZN(new_n366));
  NAND3_X1  g0166(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n365), .A2(new_n366), .B1(new_n210), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n269), .A2(new_n210), .A3(G68), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n210), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n225), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(KEYINPUT19), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n256), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n282), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n286), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n375), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n355), .A2(new_n359), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G190), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n355), .B2(new_n359), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n373), .B(new_n376), .C1(new_n223), .C2(new_n378), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n362), .A2(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n348), .A2(new_n349), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT84), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n346), .B2(new_n347), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT84), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n349), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n269), .A2(G1698), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT69), .ZN(new_n395));
  INV_X1    g0195(.A(G223), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n269), .A2(new_n298), .ZN(new_n398));
  INV_X1    g0198(.A(G222), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(new_n234), .B2(new_n269), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n292), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G45), .ZN(new_n402));
  AOI21_X1  g0202(.A(G1), .B1(new_n315), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G274), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n352), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n352), .A2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G226), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(G200), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n272), .A2(G150), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT8), .B(G58), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n370), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n256), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n285), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n217), .B1(new_n209), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(new_n217), .B2(new_n374), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT9), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n411), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT10), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n411), .A2(new_n425), .A3(new_n412), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n409), .A2(new_n339), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n421), .C1(G179), .C2(new_n409), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n295), .A2(new_n257), .ZN(new_n432));
  INV_X1    g0232(.A(G232), .ZN(new_n433));
  INV_X1    g0233(.A(G238), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n432), .B1(new_n433), .B2(new_n398), .C1(new_n395), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n292), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n407), .A2(G244), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n406), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT71), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n405), .B1(new_n435), .B2(new_n292), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(KEYINPUT71), .A3(new_n437), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n410), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(G200), .A3(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(new_n272), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n415), .B1(KEYINPUT72), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(KEYINPUT72), .B2(new_n446), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n448), .B1(new_n210), .B2(new_n234), .C1(new_n370), .C2(new_n375), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n449), .A2(new_n256), .ZN(new_n450));
  OAI21_X1  g0250(.A(G77), .B1(new_n210), .B2(G1), .ZN(new_n451));
  INV_X1    g0251(.A(new_n234), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n285), .A2(new_n451), .B1(new_n452), .B2(new_n282), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n445), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n440), .A2(new_n442), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n456), .B2(new_n305), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n440), .A2(new_n339), .A3(new_n442), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n431), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n415), .B1(new_n209), .B2(G20), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n418), .A2(new_n461), .B1(new_n374), .B2(new_n415), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n262), .A2(G33), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT7), .B(new_n210), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n202), .B1(new_n270), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G58), .A2(G68), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n203), .A2(new_n205), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n272), .A2(G159), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n284), .B1(new_n473), .B2(KEYINPUT16), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT16), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n202), .B1(new_n268), .B2(new_n270), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n472), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n463), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT17), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT76), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n259), .A2(new_n223), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G223), .A2(G1698), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n230), .B2(G1698), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n484), .B2(new_n269), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n481), .B1(new_n485), .B2(new_n291), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G41), .A2(G45), .ZN(new_n487));
  OAI21_X1  g0287(.A(G232), .B1(new_n487), .B2(G1), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n404), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n350), .B2(new_n351), .ZN(new_n490));
  OR2_X1    g0290(.A1(G223), .A2(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n230), .A2(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n264), .A2(new_n491), .A3(new_n294), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n482), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(KEYINPUT76), .A3(new_n292), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n486), .A2(new_n490), .A3(new_n410), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G200), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n310), .A2(new_n313), .B1(new_n404), .B2(new_n488), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n291), .B1(new_n493), .B2(new_n494), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT77), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n497), .A2(KEYINPUT77), .A3(new_n501), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n478), .B(new_n480), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n478), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n479), .B1(new_n506), .B2(KEYINPUT78), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n497), .A2(new_n501), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT77), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n497), .A2(KEYINPUT77), .A3(new_n501), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT79), .A4(new_n478), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n505), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n486), .A2(new_n490), .A3(new_n305), .A4(new_n496), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n339), .B1(new_n499), .B2(new_n500), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT18), .B1(new_n478), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n270), .A2(new_n466), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G68), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n470), .A2(new_n471), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT16), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n477), .A2(new_n523), .A3(new_n256), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n462), .ZN(new_n525));
  INV_X1    g0325(.A(new_n518), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT18), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n202), .A2(G20), .ZN(new_n530));
  INV_X1    g0330(.A(G77), .ZN(new_n531));
  OAI221_X1 g0331(.A(new_n530), .B1(new_n370), .B2(new_n531), .C1(new_n446), .C2(new_n217), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n256), .ZN(new_n533));
  XOR2_X1   g0333(.A(new_n533), .B(KEYINPUT11), .Z(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT73), .ZN(new_n536));
  OR3_X1    g0336(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT12), .B1(new_n282), .B2(G68), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n537), .A2(new_n538), .B1(new_n418), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n407), .A2(G238), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G97), .ZN(new_n543));
  OAI221_X1 g0343(.A(new_n543), .B1(new_n398), .B2(new_n230), .C1(new_n433), .C2(new_n394), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n292), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n545), .A3(new_n406), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(KEYINPUT13), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(KEYINPUT13), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n339), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT74), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT14), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n548), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n549), .A2(new_n553), .B1(new_n554), .B2(new_n305), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT13), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n546), .B(new_n556), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(new_n339), .A3(new_n552), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n541), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(G200), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(G190), .ZN(new_n561));
  INV_X1    g0361(.A(new_n541), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NOR4_X1   g0364(.A1(new_n460), .A2(new_n515), .A3(new_n529), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  OAI221_X1 g0366(.A(new_n566), .B1(new_n398), .B2(new_n224), .C1(new_n226), .C2(new_n394), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n292), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n314), .A2(G264), .A3(new_n320), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n305), .A3(new_n328), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n328), .A3(new_n569), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n339), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n370), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n258), .A2(G20), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n269), .A2(new_n210), .A3(G87), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT22), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g0380(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n284), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT25), .B1(new_n374), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n586), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n378), .A2(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n570), .B(new_n572), .C1(new_n585), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n584), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n583), .B1(new_n577), .B2(new_n579), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n256), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n571), .A2(G200), .ZN(new_n595));
  INV_X1    g0395(.A(new_n590), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n568), .A2(G190), .A3(new_n328), .A4(new_n569), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n300), .B(new_n210), .C1(G33), .C2(new_n225), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n256), .C1(new_n210), .C2(G116), .ZN(new_n601));
  XOR2_X1   g0401(.A(new_n601), .B(KEYINPUT20), .Z(new_n602));
  NOR2_X1   g0402(.A1(new_n282), .A2(G116), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n286), .B2(G116), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n269), .A2(G264), .A3(G1698), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI221_X1 g0407(.A(new_n606), .B1(new_n607), .B2(new_n269), .C1(new_n398), .C2(new_n226), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n292), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n314), .A2(G270), .A3(new_n320), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n328), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n611), .A3(G169), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n605), .A2(G179), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n605), .A2(new_n611), .A3(new_n616), .A4(G169), .ZN(new_n617));
  XOR2_X1   g0417(.A(KEYINPUT86), .B(KEYINPUT21), .Z(new_n618));
  AND2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(KEYINPUT85), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n605), .B1(new_n611), .B2(G200), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n410), .B2(new_n611), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n393), .A2(new_n565), .A3(new_n599), .A4(new_n625), .ZN(G372));
  NOR2_X1   g0426(.A1(new_n362), .A2(new_n380), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n598), .B1(new_n385), .B2(new_n384), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n621), .B2(new_n591), .ZN(new_n629));
  INV_X1    g0429(.A(new_n346), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n337), .A2(new_n342), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n386), .ZN(new_n633));
  XOR2_X1   g0433(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n330), .A2(new_n336), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n387), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n565), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT89), .B1(new_n519), .B2(new_n528), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n559), .A2(new_n459), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n515), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n427), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n429), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n643), .A2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n281), .A2(new_n210), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT90), .Z(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n585), .B2(new_n590), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n599), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n591), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n605), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n625), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n621), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n621), .A2(new_n662), .ZN(new_n678));
  INV_X1    g0478(.A(new_n662), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n670), .A2(new_n678), .B1(new_n667), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n213), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n365), .A2(new_n573), .A3(new_n366), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(G1), .ZN(new_n686));
  INV_X1    g0486(.A(new_n218), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  AND4_X1   g0490(.A1(new_n599), .A2(new_n621), .A3(new_n623), .A4(new_n679), .ZN(new_n691));
  AND4_X1   g0491(.A1(new_n391), .A2(new_n348), .A3(new_n349), .A4(new_n387), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n391), .B1(new_n390), .B2(new_n349), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT93), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT93), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n393), .A2(new_n696), .A3(new_n691), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n381), .A2(G179), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n568), .A2(new_n569), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n699), .A2(new_n700), .A3(new_n611), .A4(new_n338), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n381), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n338), .A3(new_n571), .A4(new_n611), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n662), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT31), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n690), .B1(new_n698), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n662), .B1(new_n631), .B2(new_n641), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n633), .A2(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n662), .B1(new_n631), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n689), .B1(new_n716), .B2(G1), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT94), .Z(G364));
  NOR2_X1   g0518(.A1(new_n280), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n209), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n683), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n674), .B2(G330), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n674), .ZN(new_n724));
  INV_X1    g0524(.A(new_n722), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n219), .B1(G20), .B2(new_n339), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n250), .A2(new_n402), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n682), .A2(new_n269), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n218), .B2(new_n402), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(new_n736), .B2(KEYINPUT95), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(KEYINPUT95), .B2(new_n736), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n682), .A2(new_n295), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n739), .A2(G355), .B1(new_n573), .B2(new_n682), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n731), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G283), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT97), .B1(new_n305), .B2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n210), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n305), .A2(KEYINPUT97), .A3(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(new_n410), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n742), .A2(new_n748), .B1(new_n750), .B2(new_n607), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(new_n305), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n410), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(G190), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G326), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G294), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n410), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n210), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(G20), .A3(new_n305), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n764), .A2(G311), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n752), .A2(G190), .A3(new_n498), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n767), .B(new_n295), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n751), .A2(new_n761), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT98), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT98), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n269), .B1(new_n769), .B2(new_n201), .ZN(new_n774));
  INV_X1    g0574(.A(new_n755), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(G159), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n202), .B1(KEYINPUT32), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n774), .B(new_n777), .C1(new_n452), .C2(new_n764), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n760), .A2(new_n225), .ZN(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n217), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(KEYINPUT32), .C2(new_n776), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n747), .A2(G107), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n749), .A2(G87), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n778), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n772), .A2(new_n773), .A3(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n725), .B(new_n741), .C1(new_n786), .C2(new_n729), .ZN(new_n787));
  INV_X1    g0587(.A(new_n728), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n674), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n724), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  INV_X1    g0591(.A(new_n454), .ZN(new_n792));
  INV_X1    g0592(.A(new_n442), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT71), .B1(new_n441), .B2(new_n437), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n305), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND4_X1   g0595(.A1(new_n792), .A2(new_n795), .A3(new_n458), .A4(new_n679), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n662), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n445), .A2(new_n454), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n443), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(new_n459), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n710), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT100), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n455), .A2(new_n797), .B1(new_n457), .B2(new_n458), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT100), .B1(new_n804), .B2(new_n796), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n801), .B1(new_n807), .B2(new_n710), .ZN(new_n808));
  INV_X1    g0608(.A(new_n709), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT101), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n722), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n729), .A2(new_n726), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n725), .B1(new_n531), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n729), .ZN(new_n816));
  INV_X1    g0616(.A(new_n769), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G143), .B1(new_n764), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  INV_X1    g0619(.A(G150), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n780), .B2(new_n819), .C1(new_n820), .C2(new_n775), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT99), .B(KEYINPUT34), .Z(new_n822));
  XNOR2_X1  g0622(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n747), .A2(G68), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n749), .A2(G50), .ZN(new_n825));
  INV_X1    g0625(.A(new_n760), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G58), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n295), .B1(new_n766), .B2(G132), .ZN(new_n828));
  AND4_X1   g0628(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n779), .B1(G283), .B2(new_n755), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n607), .B2(new_n780), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n295), .B1(new_n769), .B2(new_n758), .ZN(new_n832));
  INV_X1    g0632(.A(G311), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n763), .A2(new_n573), .B1(new_n765), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G87), .A2(new_n747), .B1(new_n749), .B2(G107), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n823), .A2(new_n829), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n815), .B1(new_n816), .B2(new_n837), .C1(new_n800), .C2(new_n727), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n813), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  INV_X1    g0640(.A(new_n277), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT35), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(KEYINPUT35), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(G116), .A3(new_n220), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT36), .Z(new_n845));
  NAND4_X1  g0645(.A1(new_n206), .A2(new_n452), .A3(G50), .A4(new_n468), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n217), .A2(G68), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n209), .B(G13), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n549), .A2(new_n553), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n552), .B1(new_n557), .B2(new_n339), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(new_n305), .C2(new_n554), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n541), .A3(new_n679), .ZN(new_n853));
  INV_X1    g0653(.A(new_n474), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n462), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n660), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n525), .B1(new_n510), .B2(new_n511), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT17), .B1(new_n859), .B2(new_n513), .ZN(new_n860));
  INV_X1    g0660(.A(new_n514), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n504), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n529), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n512), .A2(new_n513), .A3(new_n478), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n856), .B1(new_n526), .B2(new_n857), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n525), .A2(new_n526), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n525), .A2(new_n857), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n866), .A3(new_n865), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT102), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n869), .A2(KEYINPUT102), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n869), .A2(new_n874), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n858), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n515), .B2(new_n529), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n877), .A4(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n873), .A2(new_n866), .A3(new_n865), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT89), .B1(new_n478), .B2(new_n518), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT89), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n525), .A2(new_n526), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n506), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n890), .A2(new_n506), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n871), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n889), .B1(new_n897), .B2(KEYINPUT37), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n871), .B1(new_n862), .B2(new_n646), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n884), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n886), .A2(new_n887), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n865), .A2(new_n866), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n904), .A2(new_n873), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n883), .B1(new_n905), .B2(KEYINPUT102), .ZN(new_n906));
  INV_X1    g0706(.A(new_n877), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n888), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n901), .B1(new_n908), .B2(new_n884), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n884), .A2(new_n900), .A3(new_n901), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT104), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n853), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n799), .A2(new_n459), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n796), .B1(new_n710), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n541), .B(new_n662), .C1(new_n852), .C2(new_n649), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n541), .A2(new_n662), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n559), .A2(new_n563), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n884), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n646), .B2(new_n857), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n653), .B1(new_n565), .B2(new_n715), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n696), .B1(new_n393), .B2(new_n691), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n599), .A2(new_n621), .A3(new_n623), .A4(new_n679), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT93), .B(new_n927), .C1(new_n389), .C2(new_n392), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n708), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n915), .A2(new_n917), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n800), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n884), .A2(new_n900), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT40), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n698), .B2(new_n708), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT40), .B1(new_n908), .B2(new_n884), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n565), .A2(new_n929), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n690), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n925), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n209), .B2(new_n719), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n925), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n849), .B1(new_n944), .B2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n385), .A2(new_n662), .ZN(new_n947));
  MUX2_X1   g0747(.A(new_n627), .B(new_n387), .S(new_n947), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT106), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n670), .A2(new_n678), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n662), .A2(new_n288), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n630), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n637), .A2(new_n662), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n951), .A2(KEYINPUT42), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT105), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n951), .A2(new_n956), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n632), .B1(new_n956), .B2(new_n591), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(KEYINPUT42), .B1(new_n679), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n950), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n964), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n677), .A2(new_n956), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n683), .B(new_n971), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n680), .A2(new_n955), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT109), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n680), .A2(new_n955), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n676), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n670), .B2(new_n678), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n675), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(new_n951), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n716), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n987), .B2(new_n716), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n970), .B1(new_n988), .B2(new_n721), .ZN(new_n989));
  INV_X1    g0789(.A(new_n375), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n731), .B1(new_n682), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n733), .A2(new_n246), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n725), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n201), .A2(new_n750), .B1(new_n748), .B2(new_n234), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G143), .A2(new_n754), .B1(new_n755), .B2(G159), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n202), .B2(new_n760), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n764), .A2(G50), .B1(new_n766), .B2(G137), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n269), .C1(new_n820), .C2(new_n769), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n748), .A2(new_n225), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n257), .A2(new_n826), .B1(new_n754), .B2(G311), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n269), .B1(new_n766), .B2(G317), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n817), .A2(G303), .B1(new_n764), .B2(G283), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n750), .B2(new_n573), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n749), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n758), .C2(new_n775), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1000), .B(new_n1004), .C1(new_n1008), .C2(KEYINPUT111), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n999), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n993), .B1(new_n948), .B2(new_n788), .C1(new_n1012), .C2(new_n816), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n989), .A2(new_n1013), .ZN(G387));
  OAI21_X1  g0814(.A(new_n733), .B1(new_n243), .B2(new_n402), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n739), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n685), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n415), .A2(G50), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g0819(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n685), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(new_n586), .B2(new_n682), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n990), .A2(new_n826), .B1(new_n754), .B2(G159), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n415), .B2(new_n775), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n750), .A2(new_n234), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n764), .A2(G68), .B1(new_n766), .B2(G150), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1026), .B(new_n269), .C1(new_n217), .C2(new_n769), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1000), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n817), .A2(G317), .B1(new_n764), .B2(G303), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n780), .B2(new_n768), .C1(new_n833), .C2(new_n775), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n749), .A2(G294), .B1(G283), .B2(new_n826), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT49), .Z(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n269), .B1(new_n766), .B2(G326), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n748), .B2(new_n573), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1036), .B2(KEYINPUT112), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1028), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n722), .B1(new_n731), .B2(new_n1022), .C1(new_n1041), .C2(new_n816), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n671), .B2(new_n728), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n985), .B2(new_n721), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n986), .A2(new_n683), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n985), .A2(new_n716), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n981), .A2(new_n986), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n987), .A2(new_n683), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n981), .A2(new_n720), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n956), .A2(new_n728), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n731), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n225), .B2(new_n213), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n734), .A2(new_n253), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n722), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G317), .A2(new_n754), .B1(new_n817), .B2(G311), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n742), .B2(new_n750), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n775), .A2(new_n607), .B1(new_n573), .B2(new_n760), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT113), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n295), .B1(new_n765), .B2(new_n768), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G294), .B2(new_n764), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n783), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n747), .A2(G87), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n760), .A2(new_n531), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G50), .B2(new_n755), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n766), .A2(G143), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n415), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n295), .B1(new_n764), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G159), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n780), .A2(new_n820), .B1(new_n1071), .B2(new_n769), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT51), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(G68), .B2(new_n749), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1058), .A2(new_n1063), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1076), .B2(new_n729), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1050), .B1(new_n1051), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1049), .A2(new_n1078), .ZN(G390));
  OAI21_X1  g0879(.A(new_n853), .B1(new_n914), .B2(new_n918), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n903), .A2(new_n911), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n796), .B1(new_n714), .B2(new_n913), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n853), .B(new_n933), .C1(new_n1082), .C2(new_n918), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT31), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n707), .B(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n695), .B2(new_n697), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n913), .B1(new_n459), .B2(new_n662), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1087), .A2(new_n690), .A3(new_n1088), .A4(new_n918), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n929), .A2(G330), .A3(new_n800), .A4(new_n930), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1081), .A2(new_n1091), .A3(new_n1083), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n709), .A2(new_n565), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n924), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n914), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n930), .B1(new_n709), .B2(new_n800), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n1089), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1087), .A2(new_n806), .A3(new_n690), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1091), .B(new_n1082), .C1(new_n1099), .C2(new_n930), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1095), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n684), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n903), .A2(new_n911), .A3(new_n726), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n814), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n722), .B1(new_n1068), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n780), .A2(new_n742), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1065), .B(new_n1109), .C1(new_n257), .C2(new_n755), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n763), .A2(new_n225), .B1(new_n765), .B2(new_n758), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n269), .B(new_n1111), .C1(G116), .C2(new_n817), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1110), .A2(new_n1112), .A3(new_n784), .A4(new_n824), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n749), .A2(G150), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n775), .A2(new_n819), .B1(new_n780), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G159), .B2(new_n826), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n747), .A2(G50), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT114), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n764), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n766), .A2(G125), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n295), .B(new_n1123), .C1(G132), .C2(new_n817), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1113), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1108), .B1(new_n1126), .B2(new_n729), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1106), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1093), .B2(new_n720), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1105), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(G378));
  AOI22_X1  g0931(.A1(new_n755), .A2(G97), .B1(new_n764), .B2(new_n990), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT115), .Z(new_n1133));
  NOR2_X1   g0933(.A1(new_n269), .A2(G41), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n742), .B2(new_n765), .C1(new_n586), .C2(new_n769), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n780), .A2(new_n573), .B1(new_n202), .B2(new_n760), .ZN(new_n1136));
  OR3_X1    g0936(.A1(new_n1025), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1133), .B(new_n1137), .C1(G58), .C2(new_n747), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT116), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT58), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(G33), .A2(G41), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1134), .A2(G50), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1121), .A2(new_n749), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n769), .A2(new_n1116), .B1(new_n763), .B2(new_n819), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G150), .B2(new_n826), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G125), .A2(new_n754), .B1(new_n755), .B2(G132), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n766), .A2(G124), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1141), .B(new_n1149), .C1(new_n748), .C2(new_n1071), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1147), .B2(KEYINPUT59), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1140), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1139), .A2(KEYINPUT58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n729), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n725), .B1(new_n217), .B2(new_n814), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n857), .A2(new_n421), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT117), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n427), .A2(new_n429), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n427), .B2(new_n429), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1165), .A2(new_n1167), .A3(KEYINPUT118), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT118), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1155), .B(new_n1156), .C1(new_n1170), .C2(new_n727), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n939), .B2(G330), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n934), .A2(KEYINPUT40), .B1(new_n936), .B2(new_n937), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1175), .A2(new_n690), .A3(new_n1170), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n923), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1170), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n939), .A2(G330), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1173), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1175), .B2(new_n690), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n912), .C2(new_n922), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1172), .B1(new_n1183), .B2(new_n721), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1095), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1104), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1104), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n683), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1193), .A2(KEYINPUT120), .B1(new_n1186), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n1196), .A3(new_n683), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(G375));
  INV_X1    g0999(.A(new_n972), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1098), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1102), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n720), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n918), .A2(new_n726), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n722), .B1(G68), .B2(new_n1107), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1121), .A2(new_n755), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n295), .B1(new_n817), .B2(G137), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G50), .A2(new_n826), .B1(new_n754), .B2(G132), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n764), .A2(G150), .B1(new_n766), .B2(G128), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n201), .A2(new_n748), .B1(new_n750), .B2(new_n1071), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n531), .A2(new_n748), .B1(new_n750), .B2(new_n225), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n990), .A2(new_n826), .B1(new_n755), .B2(G116), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n764), .A2(new_n257), .B1(new_n766), .B2(G303), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n269), .B1(new_n817), .B2(G283), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n754), .A2(G294), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1210), .A2(new_n1211), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1205), .B1(new_n1218), .B2(new_n729), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1203), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1202), .A2(new_n1220), .ZN(G381));
  NAND4_X1  g1021(.A1(new_n989), .A2(new_n1013), .A3(new_n1049), .A4(new_n1078), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1220), .A3(new_n1202), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G378), .A2(new_n1222), .A3(new_n1225), .A4(G375), .ZN(G407));
  NOR2_X1   g1026(.A1(new_n658), .A2(G343), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT122), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1198), .A2(new_n1130), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G407), .A2(G213), .A3(new_n1229), .ZN(G409));
  XNOR2_X1  g1030(.A(new_n1201), .B(KEYINPUT60), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n683), .A3(new_n1102), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G384), .A2(new_n1220), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1220), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n839), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1237), .A2(G2897), .A3(new_n1227), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(G2897), .B2(new_n1228), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n720), .B1(new_n1183), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1177), .A2(new_n1182), .A3(KEYINPUT124), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1172), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1194), .B2(new_n972), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(KEYINPUT125), .A3(new_n1130), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1130), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1198), .B2(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1183), .A2(KEYINPUT57), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1104), .A2(new_n1189), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT119), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1104), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT120), .B1(new_n1256), .B2(new_n684), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1194), .A2(new_n1186), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1197), .A3(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(new_n1250), .A3(G378), .A4(new_n1184), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1249), .B1(new_n1251), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1228), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1240), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1265), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1259), .A2(G378), .A3(new_n1184), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT123), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1248), .B1(new_n1270), .B2(new_n1260), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(new_n1228), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1267), .B(new_n1268), .C1(new_n1272), .C2(new_n1240), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(new_n1263), .A3(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1271), .A2(new_n1227), .A3(new_n1236), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(KEYINPUT62), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1266), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1222), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(new_n790), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1281), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1222), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(KEYINPUT61), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1276), .A2(KEYINPUT63), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1237), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1271), .A2(new_n1227), .B1(new_n1239), .B2(new_n1238), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1291), .ZN(G405));
  NOR2_X1   g1092(.A1(new_n1251), .A2(new_n1261), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1198), .A2(G378), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1236), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1296), .B(new_n1285), .ZN(G402));
endmodule


