//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(new_n188), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n190), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n191), .B2(new_n195), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n197), .B2(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(G146), .B(new_n201), .C1(new_n205), .C2(new_n199), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT74), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT74), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G146), .A4(new_n201), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n198), .A2(new_n207), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n197), .A2(G110), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n201), .B1(new_n205), .B2(new_n199), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n218), .C1(new_n192), .C2(new_n193), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n221), .B(new_n223), .Z(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(new_n219), .A3(new_n224), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  AOI21_X1  g043(.A(G902), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n232), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n226), .A2(new_n234), .A3(new_n227), .A4(new_n230), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(G234), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n226), .A2(new_n227), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G472), .A2(G902), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT32), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n212), .A2(G143), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G137), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(KEYINPUT65), .A3(G137), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n269), .A3(G134), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n267), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n268), .B1(new_n267), .B2(new_n274), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n261), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n254), .A2(KEYINPUT1), .A3(new_n188), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n252), .C2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT66), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n254), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n278), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n267), .A2(new_n268), .A3(new_n274), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n263), .A2(new_n270), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n277), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G119), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n295), .A3(G116), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT69), .B1(new_n187), .B2(G116), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n190), .A2(new_n300), .A3(G116), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT2), .B(G113), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n299), .B2(new_n301), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n292), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n297), .B1(new_n190), .B2(G116), .ZN(new_n307));
  AND4_X1   g121(.A1(new_n300), .A2(new_n293), .A3(new_n295), .A4(G116), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n291), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n291), .A2(KEYINPUT30), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n277), .B(new_n315), .C1(new_n286), .C2(new_n290), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n317), .B2(new_n312), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT71), .A2(G237), .ZN(new_n322));
  AOI21_X1  g136(.A(G953), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G210), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n250), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT70), .B1(new_n309), .B2(new_n310), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n314), .B2(new_n316), .ZN(new_n332));
  INV_X1    g146(.A(new_n327), .ZN(new_n333));
  NOR4_X1   g147(.A1(new_n332), .A2(KEYINPUT31), .A3(new_n333), .A4(new_n313), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n278), .ZN(new_n338));
  INV_X1    g152(.A(new_n285), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(G128), .A3(new_n279), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n284), .B1(new_n343), .B2(new_n254), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n290), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n331), .A2(new_n347), .A3(new_n277), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n291), .A2(new_n312), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n337), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n313), .A2(KEYINPUT28), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n249), .B1(new_n335), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n315), .B1(new_n347), .B2(new_n277), .ZN(new_n354));
  INV_X1    g168(.A(new_n316), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n312), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n327), .A3(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT31), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n318), .A2(new_n250), .A3(new_n327), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n352), .A4(new_n249), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n248), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n348), .B2(new_n349), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n351), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n333), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n318), .A2(new_n333), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n327), .B1(new_n350), .B2(new_n351), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n371), .B2(KEYINPUT29), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G472), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n362), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n358), .A2(new_n352), .A3(new_n359), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n360), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT32), .B1(new_n377), .B2(new_n245), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n244), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G122), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n383), .A2(new_n386), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n305), .B2(new_n311), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n299), .B2(new_n301), .ZN(new_n398));
  OAI21_X1  g212(.A(G113), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n309), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n385), .A3(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT76), .B1(new_n382), .B2(G107), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n385), .A2(G104), .ZN(new_n404));
  OAI211_X1 g218(.A(G101), .B(new_n402), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n391), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n391), .A3(KEYINPUT77), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n381), .B1(new_n396), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n395), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n329), .B2(new_n330), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n408), .A2(new_n409), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT5), .B1(new_n307), .B2(new_n308), .ZN(new_n416));
  INV_X1    g230(.A(new_n399), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n304), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n419), .A3(new_n380), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n420), .A3(KEYINPUT6), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n261), .A2(new_n203), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n286), .B2(new_n203), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n222), .A2(G224), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n414), .A2(new_n419), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n380), .A2(KEYINPUT6), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n428), .ZN(new_n430));
  AOI211_X1 g244(.A(KEYINPUT82), .B(new_n430), .C1(new_n414), .C2(new_n419), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n421), .B(new_n425), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n396), .A2(new_n411), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT82), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n426), .A3(new_n428), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n425), .A4(new_n421), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n203), .B(new_n338), .C1(new_n339), .C2(new_n344), .ZN(new_n441));
  INV_X1    g255(.A(new_n422), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n441), .A2(new_n442), .B1(KEYINPUT7), .B2(new_n424), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n434), .B2(new_n380), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT7), .A4(new_n424), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n423), .A2(KEYINPUT86), .A3(KEYINPUT7), .A4(new_n424), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n406), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT85), .B1(new_n418), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n418), .A2(KEYINPUT84), .A3(new_n450), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n400), .B2(new_n406), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n400), .A2(new_n455), .A3(new_n406), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n451), .A2(new_n452), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n380), .B(KEYINPUT8), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n237), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n440), .A2(new_n465), .A3(new_n462), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n461), .B1(new_n433), .B2(new_n439), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT87), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  INV_X1    g286(.A(G227), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT10), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n340), .A2(G128), .B1(new_n251), .B2(new_n253), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n278), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n479), .B2(new_n406), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n261), .A2(new_n392), .A3(new_n394), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n408), .A2(KEYINPUT10), .A3(new_n409), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n480), .B(new_n481), .C1(new_n286), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n275), .A2(new_n276), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT78), .B(new_n476), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n485), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n476), .B1(new_n483), .B2(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n479), .A2(new_n406), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n345), .B2(new_n450), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT12), .A3(new_n485), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n493), .B1(new_n286), .B2(new_n406), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n345), .A2(new_n415), .A3(KEYINPUT10), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n484), .A3(new_n480), .A4(new_n481), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n476), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n237), .B1(new_n492), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n489), .A2(KEYINPUT80), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n506), .A3(new_n476), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n507), .A3(new_n500), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n476), .B1(new_n502), .B2(new_n487), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT79), .B(G469), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n504), .A2(G469), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  XOR2_X1   g328(.A(G113), .B(G122), .Z(new_n515));
  XOR2_X1   g329(.A(KEYINPUT94), .B(G104), .Z(new_n516));
  XOR2_X1   g330(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n321), .A2(new_n322), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G214), .A3(new_n222), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT89), .B1(new_n520), .B2(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(KEYINPUT89), .B2(G143), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(G214), .A3(new_n323), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n522), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT90), .B1(new_n208), .B2(new_n212), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n212), .B2(new_n208), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n205), .A2(KEYINPUT90), .A3(G146), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n524), .A3(new_n268), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n268), .B1(new_n522), .B2(new_n524), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT17), .ZN(new_n538));
  INV_X1    g352(.A(new_n218), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n522), .A2(new_n524), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n517), .B(new_n534), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n207), .A2(new_n211), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n208), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n208), .B1(KEYINPUT92), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT93), .B1(new_n550), .B2(G146), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n547), .A2(new_n552), .A3(new_n212), .A4(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n545), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n541), .A2(new_n535), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n532), .A2(new_n533), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n528), .B2(new_n526), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n554), .A2(new_n555), .B1(new_n557), .B2(new_n530), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n544), .B1(new_n558), .B2(new_n517), .ZN(new_n559));
  NOR2_X1   g373(.A1(G475), .A2(G902), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n514), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n514), .A3(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n222), .A2(G952), .ZN(new_n565));
  INV_X1    g379(.A(G234), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n320), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n237), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n252), .A2(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n188), .A2(G143), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT97), .ZN(new_n578));
  AOI21_X1  g392(.A(G134), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G116), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n580), .A2(G116), .ZN(new_n583));
  OAI21_X1  g397(.A(G107), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n385), .A3(new_n581), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n579), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n252), .A2(KEYINPUT13), .A3(G128), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n573), .B2(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT95), .B(KEYINPUT13), .C1(new_n252), .C2(G128), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n574), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n593), .A2(new_n594), .A3(G134), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n593), .B2(G134), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n587), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT14), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n583), .B1(new_n598), .B2(new_n581), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n385), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT98), .B1(new_n585), .B2(KEYINPUT14), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n577), .A2(G134), .A3(new_n578), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n603), .B(new_n586), .C1(new_n579), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT9), .B(G234), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(new_n236), .A3(G953), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n597), .A2(new_n605), .A3(new_n608), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G478), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n612), .B(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n544), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n218), .B1(new_n537), .B2(KEYINPUT17), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n555), .B2(KEYINPUT17), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n517), .B1(new_n618), .B2(new_n534), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n237), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G475), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n564), .A2(new_n572), .A3(new_n615), .A4(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G221), .B1(new_n607), .B2(G902), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n513), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G214), .B1(G237), .B2(G902), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT81), .Z(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n471), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n379), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n390), .ZN(G3));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n468), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n463), .A2(new_n466), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n469), .A2(KEYINPUT99), .A3(new_n465), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n627), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n559), .A2(new_n514), .A3(new_n560), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n621), .B1(new_n639), .B2(new_n561), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n613), .A2(new_n237), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n612), .B2(new_n613), .ZN(new_n643));
  INV_X1    g457(.A(new_n611), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n608), .B1(new_n597), .B2(new_n605), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT33), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n610), .A2(new_n647), .A3(new_n611), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(G478), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n638), .A2(new_n572), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT12), .B1(new_n495), .B2(new_n485), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n498), .A2(new_n497), .A3(new_n484), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n502), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n491), .A2(new_n488), .B1(new_n655), .B2(new_n475), .ZN(new_n656));
  OAI21_X1  g470(.A(G469), .B1(new_n656), .B2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n511), .A2(new_n512), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n624), .B(new_n243), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n377), .A2(new_n245), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n376), .B2(new_n360), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n652), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT34), .B(G104), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NOR2_X1   g480(.A1(new_n640), .A2(new_n615), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n572), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n627), .B(new_n668), .C1(new_n635), .C2(new_n637), .ZN(new_n669));
  INV_X1    g483(.A(new_n663), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(new_n629), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n220), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n241), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n239), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT101), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT37), .B(G110), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n568), .B1(new_n569), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n667), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n638), .A2(KEYINPUT102), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n469), .B2(new_n465), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n469), .A2(new_n465), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n628), .B(new_n690), .C1(new_n694), .C2(new_n636), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n624), .B1(new_n657), .B2(new_n658), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n660), .A2(new_n247), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n377), .A2(new_n248), .B1(G472), .B2(new_n372), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n680), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n691), .A2(new_n697), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(new_n318), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n327), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n348), .A2(new_n349), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n708), .B2(new_n333), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n661), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n377), .B2(new_n248), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n699), .A2(new_n704), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n704), .B1(new_n699), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n471), .B(KEYINPUT38), .Z(new_n715));
  XOR2_X1   g529(.A(new_n687), .B(KEYINPUT39), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n698), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(KEYINPUT40), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n612), .B(new_n614), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n640), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n627), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n680), .A3(new_n722), .ZN(new_n723));
  OR4_X1    g537(.A1(new_n714), .A2(new_n715), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  INV_X1    g539(.A(new_n651), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n627), .B(new_n726), .C1(new_n635), .C2(new_n637), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n701), .A3(new_n698), .A4(new_n688), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  AOI22_X1  g544(.A1(KEYINPUT80), .A2(new_n489), .B1(new_n496), .B2(new_n499), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n509), .B1(new_n731), .B2(new_n507), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n508), .A2(new_n510), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT104), .A3(new_n237), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(G469), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n623), .A3(new_n658), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n244), .B(new_n737), .C1(new_n374), .C2(new_n378), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n652), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT41), .B(G113), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  INV_X1    g555(.A(new_n668), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n638), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT105), .B1(new_n743), .B2(new_n738), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n243), .B1(new_n699), .B2(new_n700), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n669), .A2(new_n745), .A3(new_n746), .A4(new_n737), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NAND3_X1  g563(.A1(new_n736), .A2(new_n623), .A3(new_n658), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n627), .B(new_n750), .C1(new_n635), .C2(new_n637), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  INV_X1    g566(.A(new_n622), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n701), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n680), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n753), .B(new_n755), .C1(new_n374), .C2(new_n378), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n737), .B(new_n628), .C1(new_n694), .C2(new_n636), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND2_X1  g574(.A1(new_n635), .A2(new_n637), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n721), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n640), .A2(new_n720), .A3(KEYINPUT110), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n572), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n628), .A3(new_n737), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n365), .A2(KEYINPUT107), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n364), .B2(new_n351), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n333), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n246), .B1(new_n335), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT108), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n377), .A2(new_n237), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT109), .B(G472), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n776), .A3(new_n244), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n580), .ZN(G24));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n776), .A3(new_n755), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n651), .A2(new_n688), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n757), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n203), .ZN(G27));
  INV_X1    g597(.A(new_n781), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n467), .A2(new_n470), .A3(new_n628), .A4(new_n468), .ZN(new_n785));
  INV_X1    g599(.A(new_n698), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n745), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT42), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n785), .A2(new_n781), .A3(new_n786), .A4(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n378), .A2(KEYINPUT111), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n246), .B1(new_n376), .B2(new_n360), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(KEYINPUT32), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n700), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n244), .A3(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n790), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT112), .B1(new_n790), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  NAND3_X1  g615(.A1(new_n745), .A2(new_n690), .A3(new_n787), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND2_X1  g617(.A1(G469), .A2(G902), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n656), .A2(KEYINPUT45), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n656), .A2(KEYINPUT45), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(G469), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n812), .A2(KEYINPUT114), .A3(KEYINPUT46), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT114), .B1(new_n812), .B2(KEYINPUT46), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n812), .A2(KEYINPUT46), .B1(new_n511), .B2(new_n512), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n623), .A3(new_n716), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n640), .A2(new_n650), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT43), .Z(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n680), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n675), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n785), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(KEYINPUT44), .A3(new_n675), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n269), .ZN(G39));
  NAND4_X1  g642(.A1(new_n699), .A2(new_n700), .A3(new_n243), .A4(new_n784), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n785), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n623), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT47), .B1(new_n816), .B2(new_n623), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  AND2_X1   g649(.A1(new_n643), .A2(new_n649), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n640), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n640), .B2(new_n836), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n838), .A2(new_n839), .A3(new_n571), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n471), .A2(new_n840), .A3(new_n628), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n379), .A2(new_n629), .B1(new_n841), .B2(new_n663), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g658(.A(KEYINPUT116), .B1(new_n841), .B2(new_n663), .C1(new_n379), .C2(new_n629), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n471), .A2(new_n628), .A3(new_n742), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n674), .A2(new_n681), .B1(new_n846), .B2(new_n670), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n652), .A2(new_n738), .B1(new_n767), .B2(new_n777), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n747), .B2(new_n744), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n759), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n466), .B(new_n461), .C1(new_n433), .C2(new_n439), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n634), .B2(KEYINPUT87), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n628), .A3(new_n467), .A4(new_n698), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n379), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT42), .B1(new_n856), .B2(new_n784), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n791), .A2(new_n244), .A3(new_n796), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n852), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n790), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n773), .A2(new_n776), .A3(new_n755), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n784), .A3(new_n787), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n785), .A2(new_n720), .A3(new_n640), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n701), .A3(new_n698), .A4(new_n688), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n864), .A3(new_n802), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n698), .B(new_n755), .C1(new_n374), .C2(new_n378), .ZN(new_n870));
  INV_X1    g684(.A(new_n695), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(KEYINPUT102), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n782), .B1(new_n872), .B2(new_n697), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n763), .A2(new_n764), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n627), .B(new_n874), .C1(new_n635), .C2(new_n637), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n786), .A2(new_n679), .A3(new_n687), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n875), .B(new_n876), .C1(new_n712), .C2(new_n713), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n728), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n861), .A2(new_n751), .A3(new_n784), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n702), .A2(new_n877), .A3(new_n728), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n868), .A2(new_n869), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n798), .A2(new_n799), .A3(new_n865), .ZN(new_n887));
  INV_X1    g701(.A(new_n652), .ZN(new_n888));
  INV_X1    g702(.A(new_n738), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n757), .A2(new_n765), .ZN(new_n890));
  INV_X1    g704(.A(new_n777), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n888), .A2(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n748), .A3(new_n759), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n883), .A2(new_n887), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT118), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n884), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n884), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n790), .A2(new_n797), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n893), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n894), .A2(new_n897), .A3(new_n865), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n850), .A2(KEYINPUT119), .A3(new_n759), .A4(new_n905), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n883), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n885), .B1(new_n868), .B2(new_n883), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n883), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n903), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n833), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n736), .A2(new_n658), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n624), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n831), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n819), .A2(new_n567), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n777), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n824), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n627), .A3(new_n715), .A4(new_n737), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT50), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n824), .A2(new_n737), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n243), .A3(new_n567), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n714), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n930), .A2(new_n641), .A3(new_n650), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n923), .A2(new_n928), .A3(new_n780), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n925), .A2(KEYINPUT51), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT51), .B1(new_n925), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n796), .A2(new_n244), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n936), .A2(new_n923), .A3(new_n928), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT48), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n930), .A2(new_n651), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n924), .A2(new_n751), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n565), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n918), .A2(new_n942), .B1(G952), .B2(G953), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n243), .A2(new_n627), .A3(new_n624), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT49), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n818), .B(new_n944), .C1(new_n920), .C2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n945), .B2(new_n920), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n714), .A2(new_n715), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(new_n222), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n902), .A2(new_n910), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(G210), .A3(G902), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n437), .A2(new_n421), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n425), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n954), .B(new_n958), .C1(new_n953), .C2(KEYINPUT122), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(G51));
  INV_X1    g777(.A(new_n903), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n913), .B2(new_n914), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(KEYINPUT123), .A3(new_n911), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n952), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n804), .B(KEYINPUT57), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n734), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n952), .A2(G902), .A3(new_n811), .A4(new_n810), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n950), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NAND4_X1  g787(.A1(new_n952), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n974));
  INV_X1    g788(.A(new_n559), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n950), .ZN(G60));
  NAND2_X1  g792(.A1(new_n646), .A2(new_n648), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n642), .B(KEYINPUT59), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n966), .A2(new_n968), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n951), .ZN(new_n984));
  INV_X1    g798(.A(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n917), .A2(new_n912), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT54), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT53), .B1(new_n868), .B2(new_n883), .ZN(new_n988));
  OAI22_X1  g802(.A1(new_n988), .A2(KEYINPUT118), .B1(new_n896), .B2(new_n884), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n989), .B2(new_n886), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n980), .B2(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n915), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n677), .ZN(new_n996));
  INV_X1    g810(.A(new_n240), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n915), .B2(new_n994), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n951), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n951), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(G66));
  INV_X1    g817(.A(G224), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n570), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT124), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n895), .B2(G953), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n956), .B1(G898), .B2(new_n222), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G69));
  OAI21_X1  g823(.A(new_n802), .B1(new_n817), .B2(new_n826), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n875), .A2(new_n796), .A3(new_n244), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n817), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n873), .A2(new_n728), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n800), .A3(new_n834), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n222), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n317), .B(new_n550), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n686), .A2(G953), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n724), .A2(new_n728), .A3(new_n873), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT125), .ZN(new_n1023));
  OR3_X1    g837(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT62), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1023), .B1(new_n1022), .B2(KEYINPUT62), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n838), .A2(new_n839), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1027), .A2(new_n667), .ZN(new_n1028));
  NOR4_X1   g842(.A1(new_n379), .A2(new_n717), .A3(new_n785), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n817), .ZN(new_n1030));
  INV_X1    g844(.A(new_n826), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n834), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n222), .A3(new_n1017), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1021), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(G953), .B1(new_n473), .B2(new_n686), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT127), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1035), .B2(new_n851), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1043), .A2(new_n327), .A3(new_n705), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n900), .A2(new_n369), .A3(new_n706), .A4(new_n1041), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1042), .B1(new_n1015), .B2(new_n851), .ZN(new_n1046));
  INV_X1    g860(.A(new_n369), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n950), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g862(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .ZN(G57));
endmodule


