//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n458), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n461), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND4_X1  g050(.A1(new_n459), .A2(new_n462), .A3(G2105), .A4(new_n463), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n464), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(new_n464), .B2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n478), .B(new_n481), .C1(new_n485), .C2(G136), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(G114), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n476), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT68), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(new_n490), .C1(new_n476), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n498), .A2(new_n469), .A3(new_n463), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n459), .A2(new_n462), .A3(new_n463), .A4(new_n498), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n501), .B2(KEYINPUT69), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n496), .A2(KEYINPUT70), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT72), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n522), .B(new_n523), .C1(new_n519), .C2(new_n518), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n520), .A2(new_n510), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G651), .B1(G50), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G166));
  NAND2_X1  g107(.A1(new_n525), .A2(G89), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n517), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n539), .B(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(G51), .B2(new_n530), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n533), .A2(new_n538), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n537), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n530), .A2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n521), .A2(new_n524), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n530), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n535), .A2(G56), .A3(new_n536), .ZN(new_n555));
  AND2_X1   g130(.A1(G68), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n530), .A2(G53), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n517), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n567), .A2(new_n568), .B1(G651), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n525), .A2(G91), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n526), .A2(new_n531), .ZN(G303));
  NAND3_X1  g151(.A1(new_n521), .A2(new_n524), .A3(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n530), .A2(G49), .ZN(new_n578));
  AOI21_X1  g153(.A(G74), .B1(new_n535), .B2(new_n536), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n545), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n517), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G48), .B2(new_n530), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n521), .A2(new_n524), .A3(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  AND2_X1   g162(.A1(new_n537), .A2(G60), .ZN(new_n588));
  AND2_X1   g163(.A1(G72), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n530), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n525), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n530), .A2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n522), .A2(G66), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n598), .A2(KEYINPUT77), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT77), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  OR3_X1    g186(.A1(G168), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT79), .B1(G168), .B2(new_n611), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n612), .B(new_n613), .C1(G868), .C2(new_n614), .ZN(G297));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(G868), .C2(new_n614), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G860), .ZN(G148));
  OR3_X1    g193(.A1(new_n607), .A2(KEYINPUT80), .A3(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT80), .B1(new_n607), .B2(G559), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n619), .A2(G868), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n611), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n477), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n489), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n484), .C2(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n489), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  INV_X1    g212(.A(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(KEYINPUT83), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(KEYINPUT83), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n634), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n658), .A2(new_n659), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n663), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  XOR2_X1   g263(.A(G1981), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT87), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n690), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n674), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n688), .A2(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n690), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n673), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(G166), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G22), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT92), .B(G1971), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n700), .B(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(new_n703), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n705), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G6), .B(G305), .S(G16), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1981), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n714), .A2(KEYINPUT34), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT34), .B1(new_n714), .B2(new_n717), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n708), .A2(G24), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G290), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1986), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n727), .A3(G131), .ZN(new_n728));
  INV_X1    g303(.A(G131), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT89), .B1(new_n484), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G107), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  INV_X1    g310(.A(G119), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n476), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G25), .B(new_n739), .S(G29), .Z(new_n740));
  OAI211_X1 g315(.A(new_n723), .B(new_n724), .C1(new_n726), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n726), .B2(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n718), .A2(new_n719), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT36), .ZN(new_n744));
  NOR2_X1   g319(.A1(G168), .A2(new_n708), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n708), .B2(G21), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G33), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n485), .A2(G139), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G127), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n470), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  NAND2_X1  g331(.A1(G103), .A2(G2104), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G2105), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n489), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n755), .A2(G2105), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n751), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n748), .B1(new_n749), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n749), .B2(new_n763), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT24), .ZN(new_n766));
  INV_X1    g341(.A(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n762), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2084), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n746), .B2(new_n747), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n559), .B2(G16), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n708), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n614), .B2(new_n708), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT30), .B(G28), .ZN(new_n781));
  OR2_X1    g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n762), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n628), .B2(new_n762), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n772), .A2(new_n775), .A3(new_n780), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n762), .A2(G32), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n477), .A2(G129), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT26), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G105), .B2(new_n466), .ZN(new_n792));
  INV_X1    g367(.A(G141), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n792), .C1(new_n484), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n788), .B1(new_n799), .B2(new_n762), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT27), .B(G1996), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n765), .A2(new_n787), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n762), .A2(G26), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT28), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n485), .A2(G140), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(G116), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G2105), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n477), .B2(G128), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(G29), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n708), .A2(G5), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G171), .B2(new_n708), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1961), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n815), .B(new_n818), .C1(G1341), .C2(new_n774), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G4), .A2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT94), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n607), .B2(new_n708), .ZN(new_n823));
  INV_X1    g398(.A(G1348), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n762), .A2(G35), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G162), .B2(new_n762), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT29), .Z(new_n828));
  INV_X1    g403(.A(G2090), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(new_n800), .B2(new_n802), .ZN(new_n830));
  NOR2_X1   g405(.A1(G27), .A2(G29), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G164), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT98), .B(G2078), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n830), .B(new_n834), .C1(new_n829), .C2(new_n828), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n820), .A2(new_n825), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n744), .A2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n744), .A2(new_n836), .ZN(G150));
  NOR2_X1   g413(.A1(new_n607), .A2(new_n617), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n537), .A2(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n545), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n530), .A2(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n550), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n558), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n843), .A2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n559), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n840), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  AND2_X1   g433(.A1(new_n794), .A2(new_n795), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n794), .A2(new_n795), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n812), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n807), .A2(new_n811), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n796), .A2(new_n862), .A3(new_n797), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n489), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n476), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n485), .B2(G142), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(new_n863), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n861), .B2(new_n863), .ZN(new_n872));
  INV_X1    g447(.A(new_n632), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n731), .B2(new_n738), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n739), .A2(new_n632), .ZN(new_n875));
  OAI22_X1  g450(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n861), .A2(new_n863), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n868), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n870), .ZN(new_n880));
  INV_X1    g455(.A(new_n492), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n504), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n876), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n876), .B2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n761), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n880), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n761), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n876), .A2(new_n880), .A3(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n628), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n885), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n885), .A2(new_n891), .A3(KEYINPUT99), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n893), .B1(new_n885), .B2(new_n891), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(G37), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  XOR2_X1   g478(.A(G290), .B(G305), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n710), .B(G303), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n619), .A2(new_n620), .A3(new_n851), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n851), .B1(new_n619), .B2(new_n620), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n607), .A2(G299), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n596), .B(new_n614), .C1(new_n605), .C2(new_n606), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n914), .B2(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n912), .A2(KEYINPUT100), .A3(new_n916), .A4(new_n913), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n914), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n908), .B2(new_n909), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n907), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n907), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n849), .ZN(G331));
  XOR2_X1   g504(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n848), .A2(new_n850), .ZN(new_n933));
  NAND2_X1  g508(.A1(G171), .A2(G168), .ZN(new_n934));
  OAI21_X1  g509(.A(G286), .B1(new_n548), .B2(new_n552), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n851), .A2(new_n938), .A3(KEYINPUT104), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n933), .A2(new_n936), .A3(KEYINPUT103), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT103), .B1(new_n933), .B2(new_n936), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n937), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n851), .A2(new_n938), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n933), .A2(new_n936), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n921), .A2(new_n942), .B1(new_n923), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n906), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n946), .B2(new_n906), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n931), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(new_n906), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n918), .B1(new_n943), .B2(new_n944), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n914), .B1(new_n942), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n945), .A2(new_n916), .A3(new_n923), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n947), .A2(new_n957), .A3(new_n949), .A4(new_n930), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n951), .A2(new_n952), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n947), .A2(new_n957), .A3(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n946), .A2(new_n906), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(new_n949), .A3(new_n947), .A4(new_n930), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n952), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n959), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n882), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n467), .A2(G40), .A3(new_n473), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n798), .A2(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n812), .B(new_n814), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT106), .Z(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n979), .B2(new_n799), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n739), .B(new_n726), .Z(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n972), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT105), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(G1986), .B2(G290), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n972), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT110), .B1(G305), .B2(G1981), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n585), .A2(new_n586), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G305), .A2(G1981), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT107), .B(G8), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n504), .B2(new_n881), .ZN(new_n999));
  INV_X1    g574(.A(new_n970), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n988), .B(new_n710), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n1004), .B2(new_n993), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1001), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n993), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n999), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n496), .A2(KEYINPUT70), .A3(new_n504), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT70), .B1(new_n496), .B2(new_n504), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(G1384), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1000), .B(new_n1011), .C1(new_n1014), .C2(new_n1009), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1000), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n507), .A2(new_n966), .A3(new_n508), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n968), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1015), .A2(G2090), .B1(new_n1019), .B2(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT55), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n535), .A2(new_n536), .ZN(new_n1026));
  INV_X1    g601(.A(G74), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1028), .A2(G651), .B1(G49), .B2(new_n530), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(KEYINPUT108), .A3(G1976), .A4(new_n577), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G288), .B2(new_n988), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1032), .A3(new_n1001), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1030), .A2(new_n1032), .A3(new_n1036), .A4(new_n1001), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1007), .A2(new_n1008), .B1(new_n1025), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n507), .A2(new_n1009), .A3(new_n966), .A4(new_n508), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n970), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n779), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n970), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT56), .B(G2072), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1047), .C1(new_n1014), .C2(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G299), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1041), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g628(.A(KEYINPUT119), .B(new_n1051), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT115), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1019), .A2(new_n1047), .B1(new_n1044), .B2(new_n779), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT61), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n1057), .B2(new_n1051), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1057), .B2(new_n1051), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1049), .A2(KEYINPUT117), .A3(new_n1052), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n976), .B(new_n1046), .C1(new_n1014), .C2(KEYINPUT45), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n967), .B2(new_n970), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT116), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT58), .B(G1341), .Z(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT59), .B1(new_n1074), .B2(new_n559), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1076), .B(new_n558), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1067), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G2067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1015), .B2(new_n824), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n608), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1061), .A2(new_n1079), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1010), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1348), .B1(new_n1088), .B2(new_n1000), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n608), .B1(new_n1089), .B2(new_n1080), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1063), .A2(new_n1066), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1060), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT118), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1060), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n970), .A2(G2084), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1100), .B(new_n1010), .C1(new_n1018), .C2(KEYINPUT50), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n966), .A4(new_n508), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n970), .B1(new_n967), .B2(new_n968), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1966), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1088), .A2(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n747), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1110), .A3(G8), .ZN(new_n1111));
  INV_X1    g686(.A(new_n998), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G286), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1098), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1115), .A2(new_n1098), .A3(new_n1113), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1114), .A2(new_n1116), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1019), .A2(G1971), .B1(new_n1044), .B2(G2090), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1112), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1022), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1039), .A2(new_n1121), .A3(new_n1024), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(G2078), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1019), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT121), .B(G1961), .Z(new_n1127));
  AOI22_X1  g702(.A1(new_n1125), .A2(new_n1126), .B1(new_n1015), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  OAI21_X1  g704(.A(G2105), .B1(new_n472), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1129), .B2(new_n472), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n467), .A2(G40), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT123), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT124), .B(G2078), .Z(new_n1134));
  NOR3_X1   g709(.A1(new_n1133), .A2(new_n1126), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1016), .A3(new_n969), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1123), .B1(new_n1138), .B2(G171), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT53), .A4(new_n1124), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(G301), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1122), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT125), .B1(new_n1138), .B2(G171), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1128), .A2(new_n1144), .A3(G301), .A4(new_n1137), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1128), .A2(new_n1140), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1118), .B(new_n1142), .C1(new_n1148), .C2(KEYINPUT54), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1040), .B1(new_n1097), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  OAI221_X1 g727(.A(new_n1152), .B1(new_n1117), .B2(new_n1113), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1122), .A2(new_n1147), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1023), .B1(new_n1020), .B2(G8), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NOR4_X1   g732(.A1(new_n1156), .A2(new_n1115), .A3(new_n1157), .A4(G286), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT114), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1024), .A4(new_n1039), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1115), .A2(G286), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1020), .A2(G8), .ZN(new_n1162));
  OAI211_X1 g737(.A(KEYINPUT63), .B(new_n1161), .C1(new_n1162), .C2(new_n1023), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1039), .A2(new_n1024), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT114), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1039), .A2(new_n1161), .A3(new_n1121), .A4(new_n1024), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(KEYINPUT113), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1157), .B1(new_n1166), .B2(KEYINPUT113), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1160), .B(new_n1165), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n987), .B1(new_n1150), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n974), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n971), .B1(new_n1172), .B2(new_n798), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n978), .A2(KEYINPUT46), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n978), .A2(KEYINPUT46), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n739), .A2(new_n726), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n980), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n812), .A2(G2067), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n971), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n984), .A2(new_n971), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT48), .Z(new_n1183));
  OR2_X1    g758(.A1(new_n982), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1177), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g761(.A(G319), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G227), .A2(new_n1188), .ZN(new_n1189));
  AND2_X1   g763(.A1(new_n654), .A2(new_n655), .ZN(new_n1190));
  OAI211_X1 g764(.A(KEYINPUT126), .B(new_n1189), .C1(new_n1190), .C2(new_n652), .ZN(new_n1191));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1192));
  INV_X1    g766(.A(new_n1189), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1192), .B1(G401), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n697), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n697), .A2(new_n1191), .A3(KEYINPUT127), .A4(new_n1194), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n898), .A2(new_n900), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n958), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(G308));
  NAND3_X1  g776(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(G225));
endmodule


