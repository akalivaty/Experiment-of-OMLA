//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT66), .B(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n210), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n208), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AND4_X1   g0033(.A1(new_n221), .A2(new_n225), .A3(new_n226), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G222), .A2(G1698), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT69), .B(G223), .Z(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G1698), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n261), .B2(new_n256), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT68), .B(G1), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n251), .B2(new_n252), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(G226), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(G13), .A4(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G50), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n283), .A2(new_n284), .A3(new_n231), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n283), .B2(new_n231), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n264), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G50), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n201), .A2(new_n208), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G58), .ZN(new_n295));
  INV_X1    g0095(.A(G58), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT8), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(KEYINPUT71), .A3(G58), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n208), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n208), .A2(KEYINPUT72), .A3(G33), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n293), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n282), .B(new_n289), .C1(new_n307), .C2(new_n287), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n262), .A2(new_n272), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n275), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n283), .A2(new_n231), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n313), .A2(new_n291), .B1(new_n208), .B2(new_n257), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n302), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n264), .A2(new_n319), .A3(G13), .A4(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(new_n257), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(new_n312), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(G77), .A3(new_n288), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G232), .A2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G1698), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G238), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n263), .C1(G107), .C2(new_n330), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n270), .A2(new_n271), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n268), .A2(G244), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n274), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n335), .A2(new_n337), .A3(new_n309), .A4(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n327), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(G200), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n335), .A2(new_n337), .A3(G190), .A4(new_n336), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(new_n326), .A3(new_n323), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n273), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n262), .A2(new_n272), .A3(KEYINPUT74), .A4(G190), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n308), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT9), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n308), .A2(new_n353), .B1(new_n273), .B2(G200), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT10), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT10), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n350), .A2(new_n352), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n311), .B(new_n345), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n256), .B2(new_n208), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n329), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n211), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(KEYINPUT66), .A2(G68), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT66), .A2(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(G58), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n228), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT79), .ZN(new_n368));
  INV_X1    g0168(.A(G159), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n291), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G20), .A2(G33), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT79), .A3(G159), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n367), .A2(G20), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n325), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n360), .B2(new_n362), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n373), .A3(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n299), .A2(new_n300), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n287), .B2(new_n288), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n379), .A2(new_n279), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT80), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n283), .A2(new_n284), .A3(new_n231), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n264), .A2(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n301), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT80), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n379), .A2(new_n279), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n376), .A2(new_n378), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(G223), .A2(G1698), .ZN(new_n392));
  INV_X1    g0192(.A(G226), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n392), .B(new_n394), .C1(new_n254), .C2(new_n255), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n263), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n267), .A2(new_n276), .A3(new_n278), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(G232), .A3(new_n253), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n398), .A2(G190), .A3(new_n336), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n336), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n253), .B1(new_n395), .B2(new_n396), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n391), .A2(KEYINPUT82), .A3(KEYINPUT17), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n370), .A2(new_n372), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n227), .B1(new_n211), .B2(G58), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n208), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n328), .A2(new_n208), .A3(new_n329), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n212), .B1(new_n412), .B2(new_n361), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n375), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(new_n378), .A3(new_n312), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n382), .A2(new_n390), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n405), .A3(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n406), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n398), .A2(G179), .A3(new_n336), .A4(new_n400), .ZN(new_n422));
  OAI21_X1  g0222(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT18), .B1(new_n391), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n415), .A2(new_n416), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n424), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n421), .B1(KEYINPUT81), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT81), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n359), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n270), .A2(new_n436), .A3(new_n271), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G97), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n393), .A2(new_n332), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G232), .B2(new_n332), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(new_n256), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n435), .A2(new_n437), .B1(new_n441), .B2(new_n263), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n399), .A2(new_n253), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n399), .A2(new_n445), .A3(new_n253), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(G238), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT13), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n442), .B2(new_n447), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT14), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT14), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(G169), .C1(new_n449), .C2(new_n450), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n442), .A2(new_n447), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT13), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT77), .A4(new_n448), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(G179), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n452), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n324), .A2(G68), .A3(new_n288), .A4(new_n325), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT12), .A4(new_n212), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT12), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n279), .B2(G68), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n304), .A2(G77), .A3(new_n305), .ZN(new_n468));
  OAI221_X1 g0268(.A(new_n468), .B1(new_n208), .B2(new_n211), .C1(new_n281), .C2(new_n291), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT11), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n469), .A2(new_n470), .A3(new_n385), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n469), .B2(new_n385), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n463), .B(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G200), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n459), .B2(new_n455), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n473), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n457), .A2(new_n459), .A3(G190), .A4(new_n460), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(KEYINPUT78), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT78), .B1(new_n474), .B2(new_n479), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n434), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT19), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n208), .B1(new_n438), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G87), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n208), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n483), .B1(new_n302), .B2(new_n486), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n312), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n318), .A2(new_n320), .A3(new_n315), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n264), .A2(G33), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n287), .A2(new_n279), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(new_n315), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n213), .A2(new_n332), .ZN(new_n498));
  INV_X1    g0298(.A(G244), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G1698), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n500), .C1(new_n254), .C2(new_n255), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n253), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n270), .A2(G45), .A3(new_n264), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n276), .A2(new_n278), .A3(G45), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G250), .A3(new_n253), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n309), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n505), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n274), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n497), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n287), .A2(G87), .A3(new_n279), .A4(new_n495), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n493), .A3(new_n494), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n504), .A2(new_n347), .A3(new_n505), .A4(new_n507), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n475), .B1(new_n509), .B2(new_n503), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT85), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n515), .ZN(new_n518));
  INV_X1    g0318(.A(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n497), .A2(new_n508), .A3(new_n510), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n279), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n496), .B2(new_n486), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n487), .B1(new_n412), .B2(new_n361), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n531), .A2(new_n486), .A3(G107), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n371), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n527), .B1(new_n537), .B2(new_n312), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G250), .A2(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(KEYINPUT4), .A2(G244), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(G1698), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n330), .A2(new_n541), .B1(G33), .B2(G283), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n499), .A2(G1698), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n256), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n253), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT5), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G41), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G257), .B(new_n253), .C1(new_n506), .C2(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT5), .B(G41), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n270), .A2(new_n264), .A3(new_n553), .A4(G45), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(G169), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n552), .A2(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  INV_X1    g0358(.A(new_n541), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n256), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT4), .B1(new_n330), .B2(new_n544), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n263), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n562), .A3(G179), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n538), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n527), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n562), .A3(G190), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n533), .B1(new_n531), .B2(new_n530), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n567), .A2(new_n208), .B1(new_n257), .B2(new_n291), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n312), .B1(new_n568), .B2(new_n528), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n557), .A2(new_n562), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT83), .B1(new_n547), .B2(new_n555), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(G200), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(KEYINPUT84), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(new_n576), .A4(G200), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n564), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT88), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT87), .B1(new_n502), .B2(G20), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT87), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(new_n208), .A3(G33), .A4(G116), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n487), .A3(G20), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n485), .B1(new_n587), .B2(KEYINPUT22), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n330), .A2(new_n208), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  INV_X1    g0392(.A(new_n588), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n330), .A2(new_n593), .A3(new_n208), .A4(new_n589), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n586), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n208), .B1(new_n254), .B2(new_n255), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  OAI21_X1  g0398(.A(G87), .B1(new_n598), .B2(KEYINPUT86), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n588), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n600), .A3(new_n594), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n325), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT25), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n279), .B2(G107), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n487), .B2(new_n496), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n579), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n592), .B1(new_n591), .B2(new_n594), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n592), .A2(new_n596), .A3(new_n594), .A4(new_n600), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n312), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n608), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(KEYINPUT88), .A3(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(new_n253), .C1(new_n506), .C2(new_n551), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G250), .A2(G1698), .ZN(new_n616));
  INV_X1    g0416(.A(G257), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(G1698), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n330), .B1(G33), .B2(G294), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n615), .B(new_n554), .C1(new_n619), .C2(new_n253), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G179), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(G169), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n609), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n264), .B2(G33), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n324), .A2(new_n325), .A3(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n558), .B(new_n208), .C1(G33), .C2(new_n486), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(G20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n312), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n629), .A2(KEYINPUT20), .A3(new_n312), .A4(new_n630), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n318), .A2(new_n320), .A3(new_n626), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n628), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(G270), .B(new_n253), .C1(new_n506), .C2(new_n551), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n332), .A2(G264), .ZN(new_n639));
  NOR2_X1   g0439(.A1(G257), .A2(G1698), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n639), .A2(new_n640), .B1(new_n254), .B2(new_n255), .ZN(new_n641));
  INV_X1    g0441(.A(G303), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n328), .A2(new_n642), .A3(new_n329), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n263), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n638), .A2(new_n644), .A3(new_n554), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(G169), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n646), .A3(KEYINPUT21), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n638), .A2(new_n644), .A3(G179), .A4(new_n554), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n637), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT21), .B1(new_n637), .B2(new_n646), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n621), .A2(G190), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n620), .A2(G200), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n612), .A2(new_n613), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n637), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n638), .A2(new_n644), .A3(new_n554), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G190), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n657), .B(new_n659), .C1(new_n475), .C2(new_n658), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n625), .A2(new_n653), .A3(new_n656), .A4(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n482), .A2(new_n524), .A3(new_n578), .A4(new_n661), .ZN(G372));
  NAND2_X1  g0462(.A1(new_n356), .A2(new_n358), .ZN(new_n663));
  INV_X1    g0463(.A(new_n341), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n479), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n421), .B1(new_n665), .B2(new_n474), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n430), .ZN(new_n667));
  INV_X1    g0467(.A(new_n311), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n482), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n511), .B2(new_n516), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n520), .A2(KEYINPUT89), .A3(new_n522), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n624), .B1(new_n603), .B2(new_n608), .ZN(new_n675));
  INV_X1    g0475(.A(new_n652), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n650), .A4(new_n647), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n578), .A2(new_n674), .A3(new_n656), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n524), .A2(new_n564), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n563), .A2(new_n556), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n563), .B2(new_n556), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n683), .A3(new_n538), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n672), .A4(new_n673), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n678), .A2(new_n680), .A3(new_n522), .A4(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n669), .B1(new_n670), .B2(new_n688), .ZN(G369));
  AND2_X1   g0489(.A1(new_n208), .A2(G13), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n264), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n651), .B2(new_n652), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n625), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n696), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n609), .A2(new_n614), .A3(new_n696), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n625), .A2(new_n703), .A3(new_n656), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n612), .A2(new_n613), .B1(new_n622), .B2(new_n623), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n697), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n653), .B(new_n660), .C1(new_n657), .C2(new_n697), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n637), .B(new_n696), .C1(new_n651), .C2(new_n652), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n705), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n710), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n222), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n207), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n488), .A2(G116), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n720), .A2(new_n722), .B1(new_n230), .B2(new_n719), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n687), .A2(new_n725), .A3(new_n697), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n625), .A2(new_n653), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n578), .A3(new_n674), .A4(new_n656), .ZN(new_n728));
  INV_X1    g0528(.A(new_n538), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n563), .A2(new_n556), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n517), .B2(new_n523), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n511), .B1(new_n732), .B2(new_n685), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n684), .A2(new_n672), .A3(new_n673), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n728), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n725), .B1(new_n736), .B2(new_n697), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n726), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n509), .A2(new_n503), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n557), .A2(new_n562), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n620), .A4(new_n645), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n658), .A2(G179), .A3(new_n557), .A4(new_n562), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n615), .B1(new_n619), .B2(new_n253), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT93), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n502), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G238), .A2(G1698), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n499), .B2(G1698), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(new_n751), .B2(new_n330), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n505), .B(new_n507), .C1(new_n752), .C2(new_n253), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT93), .B1(new_n753), .B2(new_n745), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n744), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT30), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT94), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n742), .A2(new_n648), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n747), .B1(new_n746), .B2(new_n740), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n753), .A2(new_n745), .A3(KEYINPUT93), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n743), .B(new_n756), .C1(new_n759), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n696), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n574), .A2(KEYINPUT84), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n538), .A3(new_n577), .A4(new_n566), .ZN(new_n769));
  AND4_X1   g0569(.A1(new_n524), .A2(new_n731), .A3(new_n769), .A4(new_n697), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n770), .B2(new_n661), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(KEYINPUT95), .B(new_n743), .C1(new_n759), .C2(new_n764), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n756), .ZN(new_n775));
  AOI21_X1  g0575(.A(KEYINPUT30), .B1(new_n763), .B2(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n755), .A2(new_n758), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(KEYINPUT95), .B1(new_n778), .B2(new_n743), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n773), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n739), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n738), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n724), .B1(new_n782), .B2(G1), .ZN(G364));
  AOI21_X1  g0583(.A(new_n207), .B1(new_n690), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n719), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n715), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G330), .B2(new_n713), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n222), .A2(new_n330), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n789), .A2(new_n205), .B1(G116), .B2(new_n222), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n246), .A2(G45), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n222), .A2(new_n256), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n266), .B2(new_n230), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n208), .B1(KEYINPUT96), .B2(new_n274), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n274), .A2(KEYINPUT96), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n231), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n786), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n208), .A2(G179), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n485), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G190), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n369), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n208), .A2(new_n309), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n347), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n309), .A2(new_n475), .A3(G190), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G20), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n814), .A2(G50), .B1(G97), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n813), .A2(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G68), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n804), .A2(new_n347), .A3(G200), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n487), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n810), .A2(new_n807), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n812), .A2(new_n808), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n812), .A2(G190), .A3(new_n475), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n330), .B1(new_n825), .B2(new_n257), .C1(new_n296), .C2(new_n826), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT97), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n256), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT33), .B(G317), .Z(new_n833));
  INV_X1    g0633(.A(new_n814), .ZN(new_n834));
  INV_X1    g0634(.A(G326), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n820), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n826), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n832), .B(new_n836), .C1(G322), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n816), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n839), .A2(new_n840), .B1(new_n805), .B2(new_n642), .ZN(new_n841));
  INV_X1    g0641(.A(new_n822), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(G283), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n809), .B(KEYINPUT98), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G329), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n829), .A2(KEYINPUT97), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n830), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n803), .B1(new_n848), .B2(new_n797), .ZN(new_n849));
  INV_X1    g0649(.A(new_n800), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n713), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n788), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G396));
  NAND2_X1  g0653(.A1(new_n327), .A2(new_n696), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n344), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n341), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n664), .A2(new_n697), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n686), .B(new_n522), .C1(new_n732), .C2(new_n685), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n769), .A2(new_n731), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n707), .A2(new_n651), .A3(new_n652), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n672), .A2(new_n656), .A3(new_n673), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n697), .B(new_n859), .C1(new_n860), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n688), .A2(new_n696), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n858), .B(KEYINPUT100), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n781), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n786), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  INV_X1    g0671(.A(new_n797), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n799), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n786), .B1(new_n873), .B2(G77), .ZN(new_n874));
  INV_X1    g0674(.A(new_n825), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n837), .A2(G143), .B1(new_n875), .B2(G159), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n820), .B2(new_n292), .C1(new_n877), .C2(new_n834), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n844), .A2(G132), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n281), .A2(new_n805), .B1(new_n822), .B2(new_n821), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n256), .B(new_n883), .C1(G58), .C2(new_n816), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n485), .A2(new_n822), .B1(new_n805), .B2(new_n487), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(G283), .B2(new_n819), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n844), .A2(G311), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n256), .B1(new_n825), .B2(new_n626), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G294), .B2(new_n837), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n814), .A2(G303), .B1(G97), .B2(new_n816), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n887), .A2(new_n888), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n874), .B1(new_n893), .B2(new_n797), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n859), .B2(new_n799), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n871), .A2(new_n895), .ZN(G384));
  NOR2_X1   g0696(.A1(new_n264), .A2(new_n690), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n387), .A2(new_n389), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n378), .A2(new_n385), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n377), .B2(new_n373), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n694), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT101), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT101), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n431), .B2(new_n433), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n427), .A2(new_n424), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n427), .A2(new_n903), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n417), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n902), .A2(new_n424), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n905), .A2(new_n417), .A3(new_n907), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n917), .B2(KEYINPUT37), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n898), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n406), .A2(new_n420), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n427), .A2(new_n428), .A3(new_n424), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n428), .B1(new_n427), .B2(new_n424), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT81), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n923), .A3(new_n433), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n908), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n914), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n919), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT31), .B1(new_n765), .B2(new_n696), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n524), .A2(new_n731), .A3(new_n769), .A4(new_n697), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n625), .A2(new_n653), .A3(new_n656), .A4(new_n660), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n743), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n776), .B2(new_n777), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n772), .B1(new_n935), .B2(new_n756), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n930), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n473), .A2(new_n696), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n474), .A2(new_n479), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n474), .B2(new_n479), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n859), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT40), .B1(new_n929), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  INV_X1    g0744(.A(new_n430), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n912), .B1(new_n945), .B2(new_n920), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n911), .A2(new_n912), .A3(new_n417), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n948), .A2(new_n914), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n898), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n944), .B1(new_n928), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n942), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT104), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n942), .A3(KEYINPUT104), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT105), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n670), .A2(new_n937), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n739), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n960), .A2(KEYINPUT106), .B1(new_n957), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT106), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n928), .A2(new_n950), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n928), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n474), .A2(new_n696), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n945), .A2(new_n903), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n939), .A2(new_n940), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n857), .B2(new_n865), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n969), .B1(new_n929), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT102), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT103), .Z(new_n975));
  OAI21_X1  g0775(.A(new_n482), .B1(new_n726), .B2(new_n737), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n669), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n897), .B1(new_n962), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n962), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(G116), .A3(new_n232), .A4(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT36), .Z(new_n984));
  NAND3_X1  g0784(.A1(new_n230), .A2(G77), .A3(new_n366), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n281), .A2(G68), .ZN(new_n986));
  AOI211_X1 g0786(.A(G13), .B(new_n264), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n980), .A2(new_n988), .ZN(G367));
  NOR2_X1   g0789(.A1(new_n697), .A2(new_n519), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n511), .ZN(new_n991));
  INV_X1    g0791(.A(new_n674), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n861), .B1(new_n729), .B2(new_n696), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(new_n1000), .B1(new_n684), .B2(new_n696), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT108), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n684), .A2(new_n696), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n998), .A2(KEYINPUT107), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n701), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n696), .B1(new_n1009), .B2(new_n731), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1001), .A2(new_n706), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT42), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n996), .B(new_n997), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n625), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n697), .B1(new_n1017), .B2(new_n564), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1011), .B(KEYINPUT42), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(new_n995), .A4(new_n994), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(new_n716), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1014), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n719), .B(KEYINPUT41), .Z(new_n1027));
  NAND3_X1  g0827(.A1(new_n1001), .A2(KEYINPUT44), .A3(new_n709), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1007), .B2(new_n710), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1032));
  NAND3_X1  g0832(.A1(new_n1007), .A2(new_n710), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(new_n1007), .B2(new_n710), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n715), .A3(new_n705), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1033), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n716), .A3(new_n1031), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n700), .A2(new_n705), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT110), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n714), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n706), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(new_n706), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1043), .B2(new_n714), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1037), .A2(new_n1040), .A3(new_n782), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1027), .B1(new_n1050), .B2(new_n782), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1025), .B(new_n1026), .C1(new_n1051), .C2(new_n785), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n801), .B1(new_n222), .B2(new_n315), .C1(new_n241), .C2(new_n792), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1054), .A2(new_n786), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n825), .A2(new_n281), .B1(new_n809), .B2(new_n877), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n256), .B(new_n1057), .C1(G150), .C2(new_n837), .ZN(new_n1058));
  INV_X1    g0858(.A(G143), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n834), .C1(new_n369), .C2(new_n820), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n839), .A2(new_n821), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n296), .B2(new_n805), .C1(new_n257), .C2(new_n822), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n814), .A2(G311), .B1(G107), .B2(new_n816), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n486), .B2(new_n822), .C1(new_n840), .C2(new_n820), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n809), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n837), .A2(G303), .B1(new_n1066), .B2(G317), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT46), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n805), .B2(new_n626), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n805), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n330), .B1(new_n875), .B2(G283), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1060), .A2(new_n1063), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1056), .B1(new_n1076), .B2(new_n872), .C1(new_n993), .C2(new_n850), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1052), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G387));
  NAND2_X1  g0880(.A1(new_n1049), .A2(new_n782), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1048), .B1(new_n781), .B2(new_n738), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n719), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n702), .A2(new_n704), .A3(new_n800), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n238), .A2(new_n266), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1085), .A2(new_n792), .B1(new_n722), .B2(new_n789), .ZN(new_n1086));
  OR3_X1    g0886(.A1(new_n313), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT50), .B1(new_n313), .B2(G50), .ZN(new_n1088));
  AOI21_X1  g0888(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n722), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1086), .A2(new_n1090), .B1(new_n487), .B2(new_n718), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n786), .B1(new_n1091), .B2(new_n802), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n826), .A2(new_n281), .B1(new_n825), .B2(new_n821), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n256), .B(new_n1093), .C1(G150), .C2(new_n1066), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n814), .A2(G159), .B1(new_n842), .B2(G97), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n315), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1070), .A2(G77), .B1(new_n1096), .B2(new_n816), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n301), .A2(new_n819), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n837), .A2(G317), .B1(new_n875), .B2(G303), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n814), .A2(G322), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n831), .C2(new_n820), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT48), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1070), .A2(G294), .B1(new_n816), .B2(G283), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT49), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n256), .B1(new_n809), .B2(new_n835), .C1(new_n626), .C2(new_n822), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT114), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1108), .A2(KEYINPUT49), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1099), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1114), .B2(new_n797), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1049), .A2(new_n785), .B1(new_n1084), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1083), .A2(new_n1116), .ZN(G393));
  INV_X1    g0917(.A(new_n1040), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n716), .B1(new_n1039), .B2(new_n1031), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1081), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1050), .A3(new_n719), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n249), .A2(new_n222), .A3(new_n256), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n801), .B1(new_n486), .B2(new_n222), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G317), .A2(new_n814), .B1(new_n837), .B2(G311), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n825), .A2(new_n840), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n330), .B(new_n1127), .C1(G322), .C2(new_n1066), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n819), .A2(G303), .B1(new_n842), .B2(G107), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1070), .A2(G283), .B1(new_n816), .B2(G116), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT116), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(KEYINPUT116), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G150), .A2(new_n814), .B1(new_n837), .B2(G159), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT51), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n330), .B1(new_n809), .B2(new_n1059), .C1(new_n313), .C2(new_n825), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n820), .A2(new_n281), .B1(new_n822), .B2(new_n485), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n839), .A2(new_n257), .B1(new_n212), .B2(new_n805), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1132), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n786), .B1(new_n1122), .B2(new_n1123), .C1(new_n1140), .C2(new_n872), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1022), .B2(new_n800), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n785), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1121), .A2(new_n1144), .ZN(G390));
  NOR3_X1   g0945(.A1(new_n937), .A2(new_n941), .A3(new_n739), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n865), .A2(new_n857), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n970), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n967), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n965), .A2(new_n966), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n963), .A2(new_n1150), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n736), .A2(new_n697), .A3(new_n856), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n970), .B1(new_n1153), .B2(new_n857), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1146), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1153), .A2(new_n857), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1150), .B(new_n963), .C1(new_n1157), .C2(new_n970), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n781), .A2(new_n859), .A3(new_n1148), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT39), .B1(new_n928), .B2(new_n950), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n925), .A2(KEYINPUT38), .A3(new_n927), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT38), .B1(new_n925), .B2(new_n927), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1163), .B2(KEYINPUT39), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n971), .A2(new_n967), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1158), .B(new_n1159), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n766), .A2(new_n767), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n933), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n936), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n482), .A2(G330), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n976), .A2(new_n1172), .A3(new_n669), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1148), .B1(new_n781), .B2(new_n859), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1147), .B1(new_n1174), .B2(new_n1146), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(G330), .A3(new_n867), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n970), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1159), .A3(new_n1157), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1173), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1167), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1156), .A3(new_n1166), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n719), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1156), .A2(new_n1166), .A3(new_n785), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n786), .B1(new_n873), .B2(new_n301), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n839), .A2(new_n369), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n820), .A2(new_n877), .B1(new_n822), .B2(new_n281), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G128), .C2(new_n814), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n805), .A2(new_n292), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT53), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n844), .A2(G125), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n330), .B1(new_n825), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G132), .B2(new_n837), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .A4(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n814), .A2(G283), .B1(new_n875), .B2(G97), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n487), .B2(new_n820), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT117), .Z(new_n1198));
  AOI211_X1 g0998(.A(new_n330), .B(new_n806), .C1(G116), .C2(new_n837), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n844), .A2(G294), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n842), .A2(G68), .B1(new_n816), .B2(G77), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1195), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1185), .B1(new_n1203), .B2(new_n797), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1164), .B2(new_n799), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1184), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1183), .A2(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n663), .A2(new_n668), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n351), .A2(new_n694), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1208), .B(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT119), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n968), .A2(new_n972), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n968), .B2(new_n972), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n956), .B(G330), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n973), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n940), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n474), .A2(new_n479), .A3(new_n938), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n858), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1171), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n944), .B1(new_n1163), .B2(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n951), .A2(new_n942), .A3(KEYINPUT104), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT104), .B1(new_n951), .B2(new_n942), .ZN(new_n1228));
  OAI211_X1 g1028(.A(G330), .B(new_n1226), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n968), .A2(new_n972), .A3(new_n1216), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1221), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1219), .A2(new_n785), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1213), .A2(new_n798), .A3(new_n1215), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n786), .B1(new_n873), .B2(G50), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n330), .A2(G41), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n315), .B2(new_n825), .C1(new_n487), .C2(new_n826), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1061), .B(new_n1236), .C1(G77), .C2(new_n1070), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n834), .A2(new_n626), .B1(new_n822), .B2(new_n296), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G97), .B2(new_n819), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n844), .A2(G283), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT58), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n281), .B1(G33), .B2(G41), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n814), .A2(G125), .ZN(new_n1244));
  INV_X1    g1044(.A(G132), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n820), .B2(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n837), .A2(G128), .B1(new_n875), .B2(G137), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n805), .B2(new_n1192), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G150), .C2(new_n816), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n842), .A2(G159), .ZN(new_n1252));
  AOI211_X1 g1052(.A(G33), .B(G41), .C1(new_n1066), .C2(G124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1242), .B1(new_n1235), .B2(new_n1243), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1256), .A2(KEYINPUT118), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n872), .B1(new_n1256), .B2(KEYINPUT118), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1234), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1233), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1232), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT120), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1173), .B(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1182), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1264), .A2(KEYINPUT57), .A3(new_n1219), .A4(new_n1231), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n719), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1221), .A2(new_n1230), .A3(new_n1229), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1229), .B1(new_n1221), .B2(new_n1230), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1269), .B2(new_n1264), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1266), .B2(new_n1270), .ZN(G375));
  NOR2_X1   g1071(.A1(new_n1179), .A2(new_n1027), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1175), .A2(new_n1178), .A3(new_n1173), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n784), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n970), .A2(new_n798), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n786), .B1(new_n873), .B2(G68), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n834), .A2(new_n840), .B1(new_n805), .B2(new_n486), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G116), .B2(new_n819), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n844), .A2(G303), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n256), .B1(new_n825), .B2(new_n487), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G283), .B2(new_n837), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n842), .A2(G77), .B1(new_n1096), .B2(new_n816), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n834), .A2(new_n1245), .B1(new_n805), .B2(new_n369), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G50), .B2(new_n816), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n844), .A2(G128), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n330), .B1(new_n825), .B2(new_n292), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G137), .B2(new_n837), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1192), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n819), .A2(new_n1290), .B1(new_n842), .B2(G58), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1284), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1277), .B1(new_n1293), .B2(new_n797), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1275), .B1(new_n1276), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1274), .A2(new_n1295), .ZN(G381));
  NAND3_X1  g1096(.A1(new_n1083), .A2(new_n852), .A3(new_n1116), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1079), .A2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1299), .A2(KEYINPUT121), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(KEYINPUT121), .ZN(new_n1301));
  INV_X1    g1101(.A(G375), .ZN(new_n1302));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1301), .A3(new_n1305), .ZN(G407));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G343), .C2(new_n1304), .ZN(G409));
  NAND2_X1  g1107(.A1(G393), .A2(G396), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT113), .B1(new_n1308), .B2(new_n1297), .ZN(new_n1309));
  OR2_X1    g1109(.A1(G390), .A2(new_n1309), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1121), .A2(new_n1144), .B1(new_n1308), .B2(new_n1297), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1078), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(G390), .A2(new_n1309), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1052), .B(new_n1077), .C1(new_n1314), .C2(new_n1311), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1183), .A2(new_n1206), .A3(new_n1232), .A4(new_n1260), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1182), .A2(new_n1263), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1219), .A2(new_n1231), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1319), .A2(new_n1320), .A3(new_n1027), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(G375), .B2(G378), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n695), .A2(G213), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n719), .B1(new_n1273), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1273), .B1(new_n1179), .B2(new_n1325), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT123), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1328), .B2(new_n1327), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1330), .A2(G384), .A3(new_n1295), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G384), .B1(new_n1330), .B2(new_n1295), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1323), .A2(KEYINPUT63), .A3(new_n1324), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1317), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1323), .A2(KEYINPUT122), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT122), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT57), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(new_n719), .A3(new_n1265), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1303), .B1(new_n1341), .B2(new_n1261), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1338), .B1(new_n1342), .B2(new_n1322), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1337), .A2(new_n1343), .A3(new_n1324), .A4(new_n1333), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1335), .B1(new_n1336), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1337), .A2(new_n1343), .A3(new_n1324), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT124), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1332), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1330), .A2(G384), .A3(new_n1295), .ZN(new_n1350));
  INV_X1    g1150(.A(G2897), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1324), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1349), .A2(new_n1350), .A3(new_n1352), .ZN(new_n1353));
  OAI22_X1  g1153(.A1(new_n1331), .A2(new_n1332), .B1(new_n1351), .B2(new_n1324), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1337), .A2(new_n1343), .A3(KEYINPUT124), .A4(new_n1324), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1348), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1345), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1355), .ZN(new_n1359));
  AND2_X1   g1159(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1316), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1323), .A2(KEYINPUT62), .A3(new_n1324), .A4(new_n1333), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1362), .B(KEYINPUT125), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT62), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1344), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1361), .B1(new_n1363), .B2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1358), .B1(new_n1366), .B2(new_n1368), .ZN(G405));
  INV_X1    g1169(.A(KEYINPUT126), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1333), .A2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT127), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT127), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1333), .A2(new_n1370), .A3(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1372), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(new_n1368), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1372), .A2(new_n1367), .A3(new_n1374), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1333), .A2(new_n1370), .ZN(new_n1378));
  NOR3_X1   g1178(.A1(new_n1305), .A2(new_n1378), .A3(new_n1342), .ZN(new_n1379));
  AND3_X1   g1179(.A1(new_n1376), .A2(new_n1377), .A3(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1379), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1380), .A2(new_n1381), .ZN(G402));
endmodule


