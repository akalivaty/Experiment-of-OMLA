

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(n310), .B(KEYINPUT33), .ZN(n311) );
  XNOR2_X1 U323 ( .A(n312), .B(n311), .ZN(n315) );
  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n396) );
  INV_X1 U325 ( .A(n357), .ZN(n322) );
  XNOR2_X1 U326 ( .A(n397), .B(n396), .ZN(n572) );
  XNOR2_X1 U327 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U328 ( .A(n325), .B(n324), .ZN(n329) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n451), .B(KEYINPUT58), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G43GAT), .B(G29GAT), .Z(n291) );
  XNOR2_X1 U333 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U335 ( .A(n292), .B(KEYINPUT73), .Z(n294) );
  XNOR2_X1 U336 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n336) );
  XOR2_X1 U338 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U339 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(G218GAT), .B(G162GAT), .Z(n418) );
  XOR2_X1 U342 ( .A(KEYINPUT84), .B(n418), .Z(n298) );
  XOR2_X1 U343 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U344 ( .A(n436), .B(G106GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n300), .B(n299), .Z(n302) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n336), .B(n303), .ZN(n307) );
  XOR2_X1 U350 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n305) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G92GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(G85GAT), .B(n306), .Z(n318) );
  XNOR2_X1 U354 ( .A(n307), .B(n318), .ZN(n542) );
  XOR2_X1 U355 ( .A(KEYINPUT32), .B(KEYINPUT81), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT31), .B(KEYINPUT83), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n312) );
  AND2_X1 U358 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  INV_X1 U359 ( .A(n315), .ZN(n313) );
  NAND2_X1 U360 ( .A1(n313), .A2(KEYINPUT82), .ZN(n317) );
  INV_X1 U361 ( .A(KEYINPUT82), .ZN(n314) );
  NAND2_X1 U362 ( .A1(n315), .A2(n314), .ZN(n316) );
  NAND2_X1 U363 ( .A1(n317), .A2(n316), .ZN(n320) );
  XNOR2_X1 U364 ( .A(G204GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XOR2_X1 U367 ( .A(G176GAT), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U368 ( .A(n444), .B(n392), .ZN(n323) );
  XNOR2_X1 U369 ( .A(G57GAT), .B(KEYINPUT76), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n321), .B(KEYINPUT13), .ZN(n357) );
  XOR2_X1 U371 ( .A(G148GAT), .B(G106GAT), .Z(n327) );
  XNOR2_X1 U372 ( .A(KEYINPUT77), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U374 ( .A(KEYINPUT78), .B(n328), .Z(n429) );
  XNOR2_X1 U375 ( .A(n329), .B(n429), .ZN(n581) );
  XNOR2_X1 U376 ( .A(n581), .B(KEYINPUT41), .ZN(n562) );
  INV_X1 U377 ( .A(n562), .ZN(n548) );
  XOR2_X1 U378 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n331) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XOR2_X1 U382 ( .A(n332), .B(n419), .Z(n338) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n334) );
  XNOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT69), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U388 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n340) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G113GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n342), .B(n341), .Z(n344) );
  XOR2_X1 U392 ( .A(G169GAT), .B(G8GAT), .Z(n393) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U394 ( .A(n393), .B(n353), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n576) );
  NAND2_X1 U396 ( .A1(n548), .A2(n576), .ZN(n345) );
  NAND2_X1 U397 ( .A1(n345), .A2(KEYINPUT46), .ZN(n349) );
  INV_X1 U398 ( .A(KEYINPUT46), .ZN(n346) );
  NAND2_X1 U399 ( .A1(n576), .A2(n346), .ZN(n347) );
  OR2_X1 U400 ( .A1(n347), .A2(n562), .ZN(n348) );
  NAND2_X1 U401 ( .A1(n349), .A2(n348), .ZN(n369) );
  INV_X1 U402 ( .A(n542), .ZN(n555) );
  XOR2_X1 U403 ( .A(G155GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G78GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U406 ( .A(n353), .B(n352), .Z(n355) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U409 ( .A(n356), .B(KEYINPUT86), .Z(n359) );
  XNOR2_X1 U410 ( .A(n357), .B(KEYINPUT12), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n367) );
  XOR2_X1 U412 ( .A(G64GAT), .B(G183GAT), .Z(n361) );
  XNOR2_X1 U413 ( .A(G71GAT), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U415 ( .A(KEYINPUT85), .B(KEYINPUT14), .Z(n363) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U418 ( .A(n365), .B(n364), .Z(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n566) );
  INV_X1 U420 ( .A(n566), .ZN(n585) );
  NOR2_X1 U421 ( .A1(n555), .A2(n585), .ZN(n368) );
  AND2_X1 U422 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n370), .B(KEYINPUT47), .ZN(n377) );
  XOR2_X1 U424 ( .A(KEYINPUT112), .B(KEYINPUT45), .Z(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT65), .B(n371), .ZN(n373) );
  XNOR2_X1 U426 ( .A(KEYINPUT36), .B(n542), .ZN(n589) );
  NOR2_X1 U427 ( .A1(n566), .A2(n589), .ZN(n372) );
  XOR2_X1 U428 ( .A(n373), .B(n372), .Z(n374) );
  NOR2_X1 U429 ( .A1(n581), .A2(n374), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n576), .B(KEYINPUT75), .ZN(n557) );
  NAND2_X1 U431 ( .A1(n375), .A2(n557), .ZN(n376) );
  NAND2_X1 U432 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U433 ( .A(KEYINPUT48), .B(n378), .ZN(n527) );
  XOR2_X1 U434 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n380) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U437 ( .A(n381), .B(KEYINPUT92), .Z(n387) );
  XOR2_X1 U438 ( .A(G183GAT), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n437) );
  XOR2_X1 U441 ( .A(G204GAT), .B(G211GAT), .Z(n385) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n428) );
  XNOR2_X1 U444 ( .A(n437), .B(n428), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U446 ( .A(G92GAT), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(G36GAT), .B(G190GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n495) );
  NAND2_X1 U452 ( .A1(n527), .A2(n495), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n399) );
  XNOR2_X1 U454 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n407) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n400), .B(G127GAT), .ZN(n441) );
  XNOR2_X1 U458 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n401), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U460 ( .A(n441), .B(n426), .ZN(n405) );
  XOR2_X1 U461 ( .A(KEYINPUT6), .B(G57GAT), .Z(n403) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n415) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XOR2_X1 U467 ( .A(G85GAT), .B(G148GAT), .Z(n409) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U470 ( .A(G29GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n573) );
  INV_X1 U474 ( .A(n573), .ZN(n515) );
  XOR2_X1 U475 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n417) );
  XNOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(n418), .Z(n421) );
  XNOR2_X1 U479 ( .A(G50GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U481 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n463) );
  NAND2_X1 U487 ( .A1(n515), .A2(n463), .ZN(n432) );
  OR2_X1 U488 ( .A1(n572), .A2(n432), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n433), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U490 ( .A(KEYINPUT87), .B(KEYINPUT64), .Z(n435) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G15GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n449) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U496 ( .A(n440), .B(G176GAT), .Z(n443) );
  XNOR2_X1 U497 ( .A(n441), .B(KEYINPUT20), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G99GAT), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X2 U502 ( .A(n449), .B(n448), .Z(n530) );
  NAND2_X1 U503 ( .A1(n450), .A2(n530), .ZN(n565) );
  NOR2_X1 U504 ( .A1(n542), .A2(n565), .ZN(n453) );
  NOR2_X1 U505 ( .A1(n557), .A2(n581), .ZN(n488) );
  XOR2_X1 U506 ( .A(n495), .B(KEYINPUT94), .Z(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(n454), .ZN(n529) );
  NOR2_X1 U508 ( .A1(n530), .A2(n529), .ZN(n456) );
  XOR2_X1 U509 ( .A(n463), .B(KEYINPUT67), .Z(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT28), .B(n455), .ZN(n532) );
  NAND2_X1 U511 ( .A1(n456), .A2(n532), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n515), .A2(n457), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT95), .ZN(n472) );
  XNOR2_X1 U514 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n462) );
  NAND2_X1 U515 ( .A1(n530), .A2(n495), .ZN(n459) );
  XNOR2_X1 U516 ( .A(KEYINPUT98), .B(n459), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n460), .A2(n463), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n469) );
  INV_X1 U519 ( .A(n529), .ZN(n467) );
  XNOR2_X1 U520 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n530), .A2(n463), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT96), .B(n466), .Z(n574) );
  NAND2_X1 U524 ( .A1(n467), .A2(n574), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n515), .A2(n470), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n485) );
  NAND2_X1 U528 ( .A1(n542), .A2(n585), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U530 ( .A1(n485), .A2(n474), .ZN(n502) );
  NAND2_X1 U531 ( .A1(n488), .A2(n502), .ZN(n481) );
  NOR2_X1 U532 ( .A1(n515), .A2(n481), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT34), .B(n475), .Z(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  INV_X1 U535 ( .A(n495), .ZN(n518) );
  NOR2_X1 U536 ( .A1(n518), .A2(n481), .ZN(n477) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  INV_X1 U538 ( .A(n530), .ZN(n520) );
  NOR2_X1 U539 ( .A1(n520), .A2(n481), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n532), .A2(n481), .ZN(n483) );
  XNOR2_X1 U544 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n585), .A2(n589), .ZN(n486) );
  NAND2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .ZN(n512) );
  NAND2_X1 U550 ( .A1(n488), .A2(n512), .ZN(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT38), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n499) );
  NAND2_X1 U554 ( .A1(n573), .A2(n499), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n530), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  INV_X1 U563 ( .A(n532), .ZN(n500) );
  NAND2_X1 U564 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  NOR2_X1 U566 ( .A1(n576), .A2(n562), .ZN(n513) );
  NAND2_X1 U567 ( .A1(n513), .A2(n502), .ZN(n508) );
  NOR2_X1 U568 ( .A1(n515), .A2(n508), .ZN(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n518), .A2(n508), .ZN(n506) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n520), .A2(n508), .ZN(n507) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n532), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT108), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n515), .A2(n523), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(KEYINPUT109), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n523), .A2(n518), .ZN(n519) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n520), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n532), .ZN(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U594 ( .A1(n527), .A2(n573), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n530), .A2(n546), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT113), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U599 ( .A1(n557), .A2(n541), .ZN(n534) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  NOR2_X1 U601 ( .A1(n562), .A2(n541), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n566), .A2(n541), .ZN(n539) );
  XOR2_X1 U608 ( .A(n540), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n544) );
  XNOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  AND2_X1 U613 ( .A1(n546), .A2(n574), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n576), .A2(n554), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U617 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n585), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n565), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n561) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n564) );
  NOR2_X1 U631 ( .A1(n562), .A2(n565), .ZN(n563) );
  XOR2_X1 U632 ( .A(n564), .B(n563), .Z(G1349GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(n569), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n580) );
  XOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .Z(n578) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n588) );
  INV_X1 U643 ( .A(n588), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n586), .A2(n576), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(n580), .B(n579), .Z(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  NAND2_X1 U648 ( .A1(n586), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

