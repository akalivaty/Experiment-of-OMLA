

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n781), .ZN(n740) );
  NAND2_X1 U552 ( .A1(G8), .A2(n781), .ZN(n813) );
  NOR2_X1 U553 ( .A1(G651), .A2(n640), .ZN(n659) );
  NOR2_X1 U554 ( .A1(n775), .A2(n774), .ZN(n777) );
  OR2_X1 U555 ( .A1(n915), .A2(n737), .ZN(n738) );
  NOR2_X1 U556 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U557 ( .A1(n750), .A2(G299), .ZN(n746) );
  AND2_X1 U558 ( .A1(n731), .A2(n730), .ZN(n737) );
  NOR2_X1 U559 ( .A1(G1966), .A2(n813), .ZN(n774) );
  BUF_X1 U560 ( .A(n581), .Z(n517) );
  NOR2_X2 U561 ( .A1(n640), .A2(n520), .ZN(n656) );
  XNOR2_X1 U562 ( .A(n525), .B(KEYINPUT64), .ZN(n526) );
  NAND2_X1 U563 ( .A1(n795), .A2(n926), .ZN(n797) );
  NOR2_X2 U564 ( .A1(G651), .A2(G543), .ZN(n658) );
  NOR2_X2 U565 ( .A1(n572), .A2(n571), .ZN(G160) );
  INV_X1 U566 ( .A(KEYINPUT27), .ZN(n741) );
  XNOR2_X1 U567 ( .A(n742), .B(n741), .ZN(n744) );
  INV_X1 U568 ( .A(KEYINPUT98), .ZN(n748) );
  XNOR2_X1 U569 ( .A(n754), .B(KEYINPUT29), .ZN(n755) );
  INV_X1 U570 ( .A(KEYINPUT103), .ZN(n776) );
  INV_X1 U571 ( .A(KEYINPUT107), .ZN(n796) );
  XNOR2_X1 U572 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U573 ( .A(KEYINPUT12), .B(KEYINPUT68), .ZN(n575) );
  XNOR2_X1 U574 ( .A(n576), .B(n575), .ZN(n577) );
  INV_X1 U575 ( .A(KEYINPUT17), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n588), .A2(n587), .ZN(n933) );
  INV_X1 U577 ( .A(G651), .ZN(n520) );
  NOR2_X1 U578 ( .A1(G543), .A2(n520), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n516), .Z(n581) );
  NAND2_X1 U580 ( .A1(G65), .A2(n517), .ZN(n519) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  NAND2_X1 U582 ( .A1(G53), .A2(n659), .ZN(n518) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n524) );
  NAND2_X1 U584 ( .A1(G91), .A2(n658), .ZN(n522) );
  NAND2_X1 U585 ( .A1(G78), .A2(n656), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  OR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(G299) );
  INV_X1 U588 ( .A(G2104), .ZN(n530) );
  NOR2_X4 U589 ( .A1(G2105), .A2(n530), .ZN(n886) );
  NAND2_X1 U590 ( .A1(G102), .A2(n886), .ZN(n529) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X2 U592 ( .A(n527), .B(n526), .ZN(n568) );
  NAND2_X1 U593 ( .A1(G138), .A2(n568), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n534) );
  AND2_X1 U595 ( .A1(n530), .A2(G2105), .ZN(n889) );
  NAND2_X1 U596 ( .A1(G126), .A2(n889), .ZN(n532) );
  AND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U598 ( .A1(G114), .A2(n890), .ZN(n531) );
  NAND2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U601 ( .A1(G90), .A2(n658), .ZN(n536) );
  NAND2_X1 U602 ( .A1(G77), .A2(n656), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(KEYINPUT67), .Z(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n543) );
  NAND2_X1 U606 ( .A1(G64), .A2(n517), .ZN(n540) );
  NAND2_X1 U607 ( .A1(G52), .A2(n659), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U609 ( .A(KEYINPUT66), .B(n541), .Z(n542) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(G301) );
  INV_X1 U611 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U612 ( .A(G2451), .B(G2427), .ZN(n553) );
  XOR2_X1 U613 ( .A(G2430), .B(G2443), .Z(n545) );
  XNOR2_X1 U614 ( .A(G2435), .B(KEYINPUT110), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n545), .B(n544), .ZN(n549) );
  XOR2_X1 U616 ( .A(G2438), .B(G2454), .Z(n547) );
  XNOR2_X1 U617 ( .A(G1348), .B(G1341), .ZN(n546) );
  XNOR2_X1 U618 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U619 ( .A(n549), .B(n548), .Z(n551) );
  XNOR2_X1 U620 ( .A(G2446), .B(KEYINPUT111), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n554) );
  AND2_X1 U623 ( .A1(n554), .A2(G14), .ZN(G401) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U625 ( .A1(G123), .A2(n889), .ZN(n555) );
  XNOR2_X1 U626 ( .A(n555), .B(KEYINPUT18), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n568), .A2(G135), .ZN(n556) );
  XNOR2_X1 U628 ( .A(n556), .B(KEYINPUT82), .ZN(n557) );
  NAND2_X1 U629 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G99), .A2(n886), .ZN(n560) );
  NAND2_X1 U631 ( .A1(G111), .A2(n890), .ZN(n559) );
  NAND2_X1 U632 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n1000) );
  XNOR2_X1 U634 ( .A(n1000), .B(G2096), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n563), .B(KEYINPUT83), .ZN(n564) );
  OR2_X1 U636 ( .A1(G2100), .A2(n564), .ZN(G156) );
  INV_X1 U637 ( .A(G120), .ZN(G236) );
  INV_X1 U638 ( .A(G69), .ZN(G235) );
  INV_X1 U639 ( .A(G108), .ZN(G238) );
  NAND2_X1 U640 ( .A1(n890), .A2(G113), .ZN(n567) );
  NAND2_X1 U641 ( .A1(G101), .A2(n886), .ZN(n565) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(n565), .Z(n566) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n889), .A2(G125), .ZN(n570) );
  NAND2_X1 U645 ( .A1(G137), .A2(n568), .ZN(n569) );
  NAND2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n836) );
  NAND2_X1 U650 ( .A1(n836), .A2(G567), .ZN(n574) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U652 ( .A1(G68), .A2(n656), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G81), .A2(n658), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U655 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n579) );
  XNOR2_X1 U656 ( .A(n580), .B(n579), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n581), .A2(G56), .ZN(n582) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n582), .Z(n583) );
  NOR2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U660 ( .A(KEYINPUT70), .B(n585), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n659), .A2(G43), .ZN(n586) );
  XOR2_X1 U662 ( .A(KEYINPUT71), .B(n586), .Z(n587) );
  INV_X1 U663 ( .A(n933), .ZN(n589) );
  XNOR2_X1 U664 ( .A(G860), .B(KEYINPUT72), .ZN(n618) );
  NAND2_X1 U665 ( .A1(n589), .A2(n618), .ZN(G153) );
  INV_X1 U666 ( .A(G868), .ZN(n677) );
  NOR2_X1 U667 ( .A1(n677), .A2(G171), .ZN(n590) );
  XNOR2_X1 U668 ( .A(n590), .B(KEYINPUT73), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G54), .A2(n659), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G79), .A2(n656), .ZN(n592) );
  NAND2_X1 U671 ( .A1(G66), .A2(n517), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n658), .A2(G92), .ZN(n593) );
  XOR2_X1 U674 ( .A(KEYINPUT74), .B(n593), .Z(n594) );
  NOR2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT15), .ZN(n915) );
  INV_X1 U678 ( .A(n915), .ZN(n622) );
  NAND2_X1 U679 ( .A1(n677), .A2(n622), .ZN(n599) );
  NAND2_X1 U680 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U681 ( .A1(G63), .A2(n517), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n659), .A2(G51), .ZN(n601) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n601), .Z(n602) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n606) );
  XOR2_X1 U685 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n604) );
  XNOR2_X1 U686 ( .A(KEYINPUT6), .B(n604), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n606), .B(n605), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n658), .A2(G89), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT4), .ZN(n609) );
  NAND2_X1 U690 ( .A1(G76), .A2(n656), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U692 ( .A(KEYINPUT5), .B(n610), .Z(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n614) );
  XOR2_X1 U694 ( .A(KEYINPUT78), .B(KEYINPUT7), .Z(n613) );
  XNOR2_X1 U695 ( .A(n614), .B(n613), .ZN(G168) );
  XNOR2_X1 U696 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(G168), .ZN(G286) );
  NAND2_X1 U698 ( .A1(G868), .A2(G286), .ZN(n617) );
  NAND2_X1 U699 ( .A1(G299), .A2(n677), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(G297) );
  INV_X1 U701 ( .A(G559), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT80), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U705 ( .A(n623), .B(KEYINPUT81), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U707 ( .A1(G868), .A2(n933), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n915), .A2(G868), .ZN(n625) );
  NOR2_X1 U709 ( .A1(G559), .A2(n625), .ZN(n626) );
  NOR2_X1 U710 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U711 ( .A1(G93), .A2(n658), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G80), .A2(n656), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G67), .A2(n517), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n676) );
  XNOR2_X1 U718 ( .A(KEYINPUT84), .B(n933), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n915), .A2(G559), .ZN(n667) );
  XNOR2_X1 U720 ( .A(n634), .B(n667), .ZN(n635) );
  NOR2_X1 U721 ( .A1(G860), .A2(n635), .ZN(n636) );
  XOR2_X1 U722 ( .A(n676), .B(n636), .Z(G145) );
  NAND2_X1 U723 ( .A1(G49), .A2(n659), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U726 ( .A1(n517), .A2(n639), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G88), .A2(n658), .ZN(n644) );
  NAND2_X1 U730 ( .A1(G75), .A2(n656), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G62), .A2(n517), .ZN(n646) );
  NAND2_X1 U733 ( .A1(G50), .A2(n659), .ZN(n645) );
  NAND2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n648), .A2(n647), .ZN(G166) );
  INV_X1 U736 ( .A(G166), .ZN(G303) );
  NAND2_X1 U737 ( .A1(G85), .A2(n658), .ZN(n650) );
  NAND2_X1 U738 ( .A1(G72), .A2(n656), .ZN(n649) );
  NAND2_X1 U739 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U740 ( .A(KEYINPUT65), .B(n651), .ZN(n655) );
  NAND2_X1 U741 ( .A1(G60), .A2(n517), .ZN(n653) );
  NAND2_X1 U742 ( .A1(G47), .A2(n659), .ZN(n652) );
  AND2_X1 U743 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U744 ( .A1(n655), .A2(n654), .ZN(G290) );
  NAND2_X1 U745 ( .A1(G73), .A2(n656), .ZN(n657) );
  XNOR2_X1 U746 ( .A(n657), .B(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U747 ( .A1(G86), .A2(n658), .ZN(n661) );
  NAND2_X1 U748 ( .A1(G48), .A2(n659), .ZN(n660) );
  NAND2_X1 U749 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U750 ( .A1(G61), .A2(n517), .ZN(n662) );
  XNOR2_X1 U751 ( .A(KEYINPUT85), .B(n662), .ZN(n663) );
  NOR2_X1 U752 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U753 ( .A1(n666), .A2(n665), .ZN(G305) );
  XOR2_X1 U754 ( .A(KEYINPUT86), .B(n667), .Z(n674) );
  XNOR2_X1 U755 ( .A(G288), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U756 ( .A(G299), .B(G303), .ZN(n668) );
  XNOR2_X1 U757 ( .A(n669), .B(n668), .ZN(n671) );
  XOR2_X1 U758 ( .A(G290), .B(n933), .Z(n670) );
  XNOR2_X1 U759 ( .A(n671), .B(n670), .ZN(n673) );
  XOR2_X1 U760 ( .A(G305), .B(n676), .Z(n672) );
  XNOR2_X1 U761 ( .A(n673), .B(n672), .ZN(n903) );
  XNOR2_X1 U762 ( .A(n674), .B(n903), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n675), .A2(G868), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U766 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XOR2_X1 U767 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U768 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U771 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G235), .A2(G236), .ZN(n684) );
  XNOR2_X1 U773 ( .A(n684), .B(KEYINPUT89), .ZN(n685) );
  NOR2_X1 U774 ( .A1(G238), .A2(n685), .ZN(n686) );
  NAND2_X1 U775 ( .A1(G57), .A2(n686), .ZN(n841) );
  NAND2_X1 U776 ( .A1(G567), .A2(n841), .ZN(n693) );
  XOR2_X1 U777 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n688) );
  NAND2_X1 U778 ( .A1(G132), .A2(G82), .ZN(n687) );
  XNOR2_X1 U779 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U780 ( .A(n689), .B(KEYINPUT87), .ZN(n690) );
  NOR2_X1 U781 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G96), .A2(n691), .ZN(n842) );
  NAND2_X1 U783 ( .A1(G2106), .A2(n842), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n860) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U786 ( .A1(n860), .A2(n694), .ZN(n838) );
  NAND2_X1 U787 ( .A1(n838), .A2(G36), .ZN(G176) );
  NOR2_X1 U788 ( .A1(G164), .A2(G1384), .ZN(n726) );
  NAND2_X1 U789 ( .A1(G160), .A2(G40), .ZN(n725) );
  NOR2_X1 U790 ( .A1(n726), .A2(n725), .ZN(n830) );
  XNOR2_X1 U791 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n705) );
  NAND2_X1 U792 ( .A1(G128), .A2(n889), .ZN(n696) );
  NAND2_X1 U793 ( .A1(G116), .A2(n890), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U795 ( .A(KEYINPUT35), .B(n697), .ZN(n703) );
  NAND2_X1 U796 ( .A1(G104), .A2(n886), .ZN(n699) );
  NAND2_X1 U797 ( .A1(G140), .A2(n568), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n701) );
  XOR2_X1 U799 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n700) );
  XNOR2_X1 U800 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U802 ( .A(n705), .B(n704), .ZN(n881) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NOR2_X1 U804 ( .A1(n881), .A2(n828), .ZN(n991) );
  NAND2_X1 U805 ( .A1(n830), .A2(n991), .ZN(n825) );
  NAND2_X1 U806 ( .A1(G129), .A2(n889), .ZN(n707) );
  NAND2_X1 U807 ( .A1(G117), .A2(n890), .ZN(n706) );
  NAND2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U809 ( .A(KEYINPUT92), .B(n708), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n886), .A2(G105), .ZN(n709) );
  XOR2_X1 U811 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U812 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U813 ( .A1(G141), .A2(n568), .ZN(n712) );
  NAND2_X1 U814 ( .A1(n713), .A2(n712), .ZN(n897) );
  NAND2_X1 U815 ( .A1(n897), .A2(G1996), .ZN(n721) );
  NAND2_X1 U816 ( .A1(G119), .A2(n889), .ZN(n715) );
  NAND2_X1 U817 ( .A1(G107), .A2(n890), .ZN(n714) );
  NAND2_X1 U818 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U819 ( .A1(G95), .A2(n886), .ZN(n717) );
  NAND2_X1 U820 ( .A1(G131), .A2(n568), .ZN(n716) );
  NAND2_X1 U821 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U822 ( .A1(n719), .A2(n718), .ZN(n877) );
  NAND2_X1 U823 ( .A1(G1991), .A2(n877), .ZN(n720) );
  NAND2_X1 U824 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U825 ( .A(n722), .B(KEYINPUT93), .ZN(n1002) );
  XOR2_X1 U826 ( .A(n830), .B(KEYINPUT94), .Z(n723) );
  NOR2_X1 U827 ( .A1(n1002), .A2(n723), .ZN(n822) );
  INV_X1 U828 ( .A(n822), .ZN(n724) );
  NAND2_X1 U829 ( .A1(n825), .A2(n724), .ZN(n817) );
  XNOR2_X1 U830 ( .A(n725), .B(KEYINPUT95), .ZN(n727) );
  NAND2_X2 U831 ( .A1(n727), .A2(n726), .ZN(n781) );
  NOR2_X1 U832 ( .A1(G2084), .A2(n781), .ZN(n761) );
  NAND2_X1 U833 ( .A1(G8), .A2(n761), .ZN(n779) );
  AND2_X1 U834 ( .A1(n781), .A2(G1341), .ZN(n728) );
  NOR2_X1 U835 ( .A1(n728), .A2(n933), .ZN(n731) );
  INV_X1 U836 ( .A(G1996), .ZN(n967) );
  NOR2_X1 U837 ( .A1(n781), .A2(n967), .ZN(n729) );
  XOR2_X1 U838 ( .A(n729), .B(KEYINPUT26), .Z(n730) );
  NAND2_X1 U839 ( .A1(n737), .A2(n915), .ZN(n736) );
  INV_X1 U840 ( .A(G2067), .ZN(n965) );
  NOR2_X1 U841 ( .A1(n781), .A2(n965), .ZN(n732) );
  XNOR2_X1 U842 ( .A(n732), .B(KEYINPUT97), .ZN(n734) );
  NAND2_X1 U843 ( .A1(n781), .A2(G1348), .ZN(n733) );
  NAND2_X1 U844 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U845 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U846 ( .A1(n739), .A2(n738), .ZN(n747) );
  NAND2_X1 U847 ( .A1(n740), .A2(G2072), .ZN(n742) );
  NAND2_X1 U848 ( .A1(G1956), .A2(n781), .ZN(n743) );
  NAND2_X1 U849 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U850 ( .A(n745), .B(KEYINPUT96), .ZN(n750) );
  NAND2_X1 U851 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U852 ( .A(n749), .B(n748), .ZN(n753) );
  NAND2_X1 U853 ( .A1(n750), .A2(G299), .ZN(n751) );
  XOR2_X1 U854 ( .A(n751), .B(KEYINPUT28), .Z(n752) );
  NOR2_X1 U855 ( .A1(n753), .A2(n752), .ZN(n756) );
  INV_X1 U856 ( .A(KEYINPUT99), .ZN(n754) );
  XNOR2_X1 U857 ( .A(n756), .B(n755), .ZN(n760) );
  INV_X1 U858 ( .A(G1961), .ZN(n938) );
  NAND2_X1 U859 ( .A1(n781), .A2(n938), .ZN(n758) );
  XNOR2_X1 U860 ( .A(KEYINPUT25), .B(G2078), .ZN(n973) );
  NAND2_X1 U861 ( .A1(n740), .A2(n973), .ZN(n757) );
  NAND2_X1 U862 ( .A1(n758), .A2(n757), .ZN(n767) );
  NAND2_X1 U863 ( .A1(G171), .A2(n767), .ZN(n759) );
  NAND2_X1 U864 ( .A1(n760), .A2(n759), .ZN(n773) );
  NOR2_X1 U865 ( .A1(n761), .A2(n774), .ZN(n762) );
  NAND2_X1 U866 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U867 ( .A(KEYINPUT101), .B(n763), .ZN(n765) );
  XOR2_X1 U868 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n764) );
  XNOR2_X1 U869 ( .A(n765), .B(n764), .ZN(n766) );
  NOR2_X1 U870 ( .A1(G168), .A2(n766), .ZN(n769) );
  NOR2_X1 U871 ( .A1(G171), .A2(n767), .ZN(n768) );
  NOR2_X1 U872 ( .A1(n769), .A2(n768), .ZN(n771) );
  XOR2_X1 U873 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n770) );
  XNOR2_X1 U874 ( .A(n771), .B(n770), .ZN(n772) );
  NAND2_X1 U875 ( .A1(n773), .A2(n772), .ZN(n780) );
  INV_X1 U876 ( .A(n780), .ZN(n775) );
  XNOR2_X1 U877 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U878 ( .A1(n779), .A2(n778), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n780), .A2(G286), .ZN(n787) );
  NOR2_X1 U880 ( .A1(G1971), .A2(n813), .ZN(n783) );
  NOR2_X1 U881 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U882 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U883 ( .A(n784), .B(KEYINPUT104), .ZN(n785) );
  NAND2_X1 U884 ( .A1(n785), .A2(G303), .ZN(n786) );
  NAND2_X1 U885 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n788), .A2(G8), .ZN(n789) );
  XNOR2_X1 U887 ( .A(n789), .B(KEYINPUT32), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n805) );
  NOR2_X1 U889 ( .A1(G1976), .A2(G288), .ZN(n800) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n800), .A2(n792), .ZN(n925) );
  XOR2_X1 U892 ( .A(n925), .B(KEYINPUT105), .Z(n793) );
  NAND2_X1 U893 ( .A1(n805), .A2(n793), .ZN(n795) );
  NAND2_X1 U894 ( .A1(G288), .A2(G1976), .ZN(n794) );
  XNOR2_X1 U895 ( .A(n794), .B(KEYINPUT106), .ZN(n926) );
  NOR2_X1 U896 ( .A1(n813), .A2(n798), .ZN(n799) );
  NOR2_X1 U897 ( .A1(KEYINPUT33), .A2(n799), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n800), .A2(KEYINPUT33), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n801), .A2(n813), .ZN(n802) );
  XOR2_X1 U900 ( .A(G1981), .B(G305), .Z(n922) );
  NAND2_X1 U901 ( .A1(n804), .A2(n922), .ZN(n810) );
  NOR2_X1 U902 ( .A1(G2090), .A2(G303), .ZN(n806) );
  NAND2_X1 U903 ( .A1(G8), .A2(n806), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n805), .A2(n807), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n808), .A2(n813), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n815) );
  NOR2_X1 U907 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U908 ( .A(n811), .B(KEYINPUT24), .Z(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n819) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U913 ( .A1(n919), .A2(n830), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n833) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n897), .ZN(n989) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n877), .ZN(n1004) );
  NOR2_X1 U918 ( .A1(n820), .A2(n1004), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n989), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT108), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n881), .A2(n828), .ZN(n993) );
  NAND2_X1 U925 ( .A1(n829), .A2(n993), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U928 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n834) );
  XNOR2_X1 U929 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G1), .A2(G3), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n840), .B(KEYINPUT112), .ZN(G188) );
  INV_X1 U937 ( .A(G132), .ZN(G219) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G82), .ZN(G220) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1961), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1981), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(G2474), .B(G1956), .Z(n857) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G229) );
  XNOR2_X1 U961 ( .A(KEYINPUT113), .B(n860), .ZN(G319) );
  NAND2_X1 U962 ( .A1(G124), .A2(n889), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n568), .A2(G136), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(KEYINPUT114), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G100), .A2(n886), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G112), .A2(n890), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G130), .A2(n889), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G118), .A2(n890), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n886), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G142), .A2(n568), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U977 ( .A(KEYINPUT115), .B(n873), .ZN(n874) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n874), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n885) );
  XNOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n877), .B(KEYINPUT116), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U984 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n899) );
  NAND2_X1 U987 ( .A1(G103), .A2(n886), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G139), .A2(n568), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G127), .A2(n889), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G115), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(KEYINPUT117), .B(n893), .ZN(n894) );
  XNOR2_X1 U994 ( .A(KEYINPUT47), .B(n894), .ZN(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n994) );
  XNOR2_X1 U996 ( .A(n897), .B(n994), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U998 ( .A(G162), .B(n1000), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(G286), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(G171), .B(n915), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n907), .Z(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT118), .B(n908), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  XOR2_X1 U1009 ( .A(KEYINPUT119), .B(n909), .Z(n910) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n911), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .ZN(n937) );
  XOR2_X1 U1016 ( .A(G1956), .B(G299), .Z(n914) );
  XNOR2_X1 U1017 ( .A(n914), .B(KEYINPUT126), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(G1348), .B(n915), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(KEYINPUT57), .B(n924), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G1961), .B(G301), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1031 ( .A(G1341), .B(n933), .Z(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n1018) );
  XNOR2_X1 U1034 ( .A(G5), .B(n938), .ZN(n956) );
  XNOR2_X1 U1035 ( .A(KEYINPUT59), .B(G4), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(KEYINPUT127), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G1348), .B(n940), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G19), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1956), .B(G20), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(KEYINPUT60), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G1986), .B(G24), .Z(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G21), .B(G1966), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT61), .B(n959), .ZN(n961) );
  INV_X1 U1056 ( .A(G16), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n962), .A2(G11), .ZN(n1016) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G25), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G26), .B(n965), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n966), .A2(G28), .ZN(n970) );
  XOR2_X1 U1064 ( .A(KEYINPUT122), .B(n967), .Z(n968) );
  XNOR2_X1 U1065 ( .A(G32), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G27), .B(n973), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1070 ( .A(n976), .B(KEYINPUT123), .Z(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n977), .ZN(n980) );
  XOR2_X1 U1072 ( .A(G35), .B(G2090), .Z(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(KEYINPUT124), .ZN(n984) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n982), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n986), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n987), .B(KEYINPUT55), .ZN(n1014) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT51), .B(n990), .Z(n1010) );
  INV_X1 U1085 ( .A(n991), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1008) );
  XOR2_X1 U1087 ( .A(G2072), .B(n994), .Z(n996) );
  XOR2_X1 U1088 ( .A(G164), .B(G2078), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT120), .B(n997), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT50), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(G2084), .B(G160), .Z(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(G29), .A2(n1012), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

