//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n642, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G173));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n459), .A2(G567), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(new_n463));
  NAND2_X1  g038(.A1(new_n457), .A2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n475), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G125), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(new_n486), .B1(G113), .B2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n479), .B1(new_n487), .B2(new_n474), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT70), .ZN(G160));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n472), .A2(new_n473), .A3(G2105), .A4(new_n475), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n476), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G136), .B2(new_n495), .ZN(G162));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n474), .A2(G114), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(new_n498), .A3(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n504), .B1(new_n492), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n473), .A2(new_n475), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n508), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n499), .A2(new_n497), .A3(new_n501), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n503), .B2(new_n498), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G138), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(G2105), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n508), .A2(KEYINPUT73), .A3(new_n472), .A4(new_n516), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n472), .A2(new_n473), .A3(new_n516), .A4(new_n475), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(KEYINPUT4), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(new_n474), .A3(G138), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n481), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n523), .A4(new_n516), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n507), .A2(new_n514), .B1(new_n521), .B2(new_n527), .ZN(G164));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT76), .A2(G651), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n530), .B(KEYINPUT6), .C1(KEYINPUT75), .C2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G50), .A2(G543), .ZN(new_n536));
  AND2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G75), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G62), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT75), .B(G651), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(G303));
  INV_X1    g123(.A(G303), .ZN(G166));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT7), .Z(new_n551));
  INV_X1    g126(.A(new_n539), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n552), .A2(G63), .A3(G651), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n534), .A2(new_n539), .ZN(new_n554));
  AOI211_X1 g129(.A(new_n551), .B(new_n553), .C1(new_n554), .C2(G89), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n534), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n532), .A2(KEYINPUT77), .A3(new_n533), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n557), .A2(G543), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G51), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n555), .A2(new_n560), .ZN(G286));
  INV_X1    g136(.A(G286), .ZN(G168));
  NAND2_X1  g137(.A1(G77), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G64), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n539), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(new_n546), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(G90), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n535), .A2(new_n552), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n559), .A2(G52), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(G171));
  NAND2_X1  g147(.A1(new_n559), .A2(G43), .ZN(new_n573));
  NAND2_X1  g148(.A1(G68), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G56), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n539), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n554), .A2(G81), .B1(new_n546), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  INV_X1    g159(.A(G91), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT79), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT80), .B(G65), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n587), .B1(new_n552), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n569), .A2(new_n585), .B1(new_n589), .B2(new_n529), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n557), .A2(G543), .A3(new_n558), .ZN(new_n591));
  INV_X1    g166(.A(G53), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT9), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n534), .B2(new_n556), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT9), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n595), .A2(new_n596), .A3(G53), .A4(new_n558), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n590), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(G299));
  INV_X1    g177(.A(G171), .ZN(G301));
  NAND3_X1  g178(.A1(new_n595), .A2(G49), .A3(new_n558), .ZN(new_n604));
  INV_X1    g179(.A(G74), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n529), .B1(new_n539), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n554), .B2(G87), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G288));
  NAND2_X1  g184(.A1(G48), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G86), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n539), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n535), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G73), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G61), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n539), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n546), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G305));
  XOR2_X1   g193(.A(KEYINPUT83), .B(G85), .Z(new_n619));
  NAND2_X1  g194(.A1(G72), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G60), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n539), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n554), .A2(new_n619), .B1(new_n546), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT82), .B(G47), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n591), .B2(new_n624), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n554), .A2(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n559), .A2(G54), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n552), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(new_n529), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n626), .B1(new_n634), .B2(G868), .ZN(G321));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NOR2_X1   g212(.A1(G286), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G299), .B(KEYINPUT85), .Z(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(new_n637), .ZN(G297));
  XNOR2_X1  g215(.A(G297), .B(KEYINPUT86), .ZN(G280));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n634), .B1(new_n642), .B2(G860), .ZN(G148));
  NAND2_X1  g218(.A1(new_n634), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G868), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n484), .A2(new_n468), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT13), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n650), .A2(new_n651), .B1(KEYINPUT87), .B2(G2100), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n495), .A2(G135), .ZN(new_n656));
  INV_X1    g231(.A(new_n492), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G123), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n474), .A2(G111), .ZN(new_n659));
  OAI21_X1  g234(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n656), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2096), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n662), .ZN(G156));
  XOR2_X1   g238(.A(KEYINPUT15), .B(G2435), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT89), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2427), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT88), .B(G2438), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT14), .ZN(new_n671));
  XOR2_X1   g246(.A(G2451), .B(G2454), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(G14), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(new_n676), .ZN(G401));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2072), .B(G2078), .Z(new_n683));
  XNOR2_X1  g258(.A(G2067), .B(G2678), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n683), .A2(KEYINPUT90), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n689), .A3(new_n685), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n683), .B(KEYINPUT17), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n682), .C1(new_n691), .C2(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n685), .A3(new_n681), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2096), .B(G2100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1971), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n701), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT20), .Z(new_n705));
  AOI211_X1 g280(.A(new_n703), .B(new_n705), .C1(new_n698), .C2(new_n702), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT99), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT26), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n495), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n657), .A2(G129), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G32), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT27), .Z(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G4), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n634), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT97), .B(G1348), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n724), .A2(G1996), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n725), .A2(G20), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT103), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT23), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT104), .B(G1956), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G168), .A2(new_n725), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n725), .B2(G21), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT101), .B(G1966), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT102), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n579), .B2(G16), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G1341), .Z(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n725), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n725), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(new_n474), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n495), .A2(G139), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G33), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n758), .A2(G2072), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(G2072), .B1(new_n758), .B2(new_n760), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT30), .B(G28), .ZN(new_n763));
  INV_X1    g338(.A(G29), .ZN(new_n764));
  OR2_X1    g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  NAND2_X1  g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n661), .B2(new_n764), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n761), .A2(new_n762), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n764), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  OR2_X1    g346(.A1(G104), .A2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n772), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n773));
  INV_X1    g348(.A(G128), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n492), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G140), .B2(new_n495), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(new_n764), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n739), .A2(new_n740), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n750), .A2(new_n769), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(KEYINPUT24), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT24), .B2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(G160), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n764), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  NOR2_X1   g362(.A1(G164), .A2(new_n764), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G27), .B2(new_n764), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n786), .A2(new_n787), .B1(new_n443), .B2(new_n789), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n742), .A2(new_n749), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n786), .A2(new_n787), .B1(new_n443), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n764), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n764), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT29), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n724), .B2(G1996), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n731), .A2(new_n737), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n725), .A2(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n608), .B2(new_n725), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n725), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n725), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n725), .A2(G6), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n613), .A2(new_n617), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n725), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT95), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n805), .A2(new_n806), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n764), .A2(G25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n657), .A2(G119), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n474), .A2(G107), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n495), .A2(KEYINPUT91), .A3(G131), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT91), .B1(new_n495), .B2(G131), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT92), .Z(new_n829));
  OAI21_X1  g404(.A(new_n822), .B1(new_n829), .B2(new_n764), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT93), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G1991), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  MUX2_X1   g410(.A(G24), .B(G290), .S(G16), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n800), .B1(new_n840), .B2(new_n841), .ZN(G311));
  INV_X1    g417(.A(new_n800), .ZN(new_n843));
  INV_X1    g418(.A(new_n841), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G150));
  XNOR2_X1  g421(.A(KEYINPUT105), .B(G55), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n559), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n539), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n554), .A2(G93), .B1(new_n546), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n634), .A2(G559), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT106), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n573), .A2(new_n848), .A3(new_n577), .A4(new_n852), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n573), .A2(new_n577), .B1(new_n848), .B2(new_n852), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n857), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n868), .B1(new_n863), .B2(new_n867), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n855), .B1(new_n871), .B2(new_n872), .ZN(G145));
  XNOR2_X1  g448(.A(G160), .B(new_n661), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n495), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n657), .A2(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n474), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n650), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n829), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n776), .B1(new_n720), .B2(new_n721), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n720), .A2(new_n721), .A3(new_n776), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n829), .B1(new_n888), .B2(new_n884), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n520), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT4), .B1(new_n518), .B2(new_n519), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n527), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n506), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n889), .A3(new_n882), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n506), .B1(new_n521), .B2(new_n527), .ZN(new_n899));
  INV_X1    g474(.A(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n901), .A3(new_n757), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n757), .B1(new_n898), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n876), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n756), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n875), .A3(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g486(.A1(new_n853), .A2(new_n637), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n644), .B(new_n862), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n633), .B1(new_n600), .B2(new_n601), .ZN(new_n914));
  INV_X1    g489(.A(new_n633), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n593), .A2(new_n597), .ZN(new_n916));
  INV_X1    g491(.A(new_n590), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT81), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n920), .A3(new_n599), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n914), .A2(new_n921), .A3(KEYINPUT41), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n913), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n914), .A2(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n913), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n608), .B(G166), .ZN(new_n928));
  XNOR2_X1  g503(.A(G290), .B(G305), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n927), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n912), .B1(new_n932), .B2(new_n637), .ZN(G295));
  OAI21_X1  g508(.A(new_n912), .B1(new_n932), .B2(new_n637), .ZN(G331));
  NAND2_X1  g509(.A1(new_n578), .A2(new_n853), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n935), .A2(G286), .A3(new_n859), .ZN(new_n936));
  AOI21_X1  g511(.A(G286), .B1(new_n935), .B2(new_n859), .ZN(new_n937));
  OAI21_X1  g512(.A(G301), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(G168), .B1(new_n860), .B2(new_n861), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(G286), .A3(new_n859), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(G171), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n942), .A2(KEYINPUT107), .A3(new_n925), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT107), .B1(new_n942), .B2(new_n925), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n941), .B(new_n938), .C1(new_n923), .C2(new_n922), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n930), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n925), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n942), .A2(KEYINPUT107), .A3(new_n925), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n947), .A3(new_n930), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT108), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n947), .A3(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(new_n930), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n948), .A2(new_n954), .A3(new_n909), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n947), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n956), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n953), .B2(KEYINPUT108), .ZN(new_n965));
  AND4_X1   g540(.A1(KEYINPUT43), .A2(new_n964), .A3(new_n965), .A4(new_n948), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n965), .A3(new_n959), .A4(new_n948), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n896), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT45), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n894), .B2(new_n895), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT111), .B(G40), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n479), .B(new_n982), .C1(new_n487), .C2(new_n474), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT112), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n776), .B(new_n778), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT113), .Z(new_n994));
  XNOR2_X1  g569(.A(new_n722), .B(G1996), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n984), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n883), .A2(new_n833), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n829), .A2(new_n832), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n984), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n985), .A2(G1996), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT46), .Z(new_n1002));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n984), .B1(new_n722), .B2(new_n992), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT125), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n991), .A2(new_n1000), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n996), .A2(new_n997), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n776), .A2(new_n778), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n985), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1956), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G113), .A2(G2104), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n485), .B1(new_n484), .B2(G125), .ZN(new_n1016));
  AND4_X1   g591(.A1(new_n485), .A2(new_n480), .A3(new_n475), .A4(G125), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n981), .B(new_n478), .C1(new_n1018), .C2(G2105), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n1020));
  OAI211_X1 g595(.A(new_n1014), .B(new_n1019), .C1(new_n978), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n510), .B1(new_n509), .B2(new_n513), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n894), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n974), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1020), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n899), .B2(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1014), .B1(new_n1029), .B2(new_n1019), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1013), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(KEYINPUT57), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(KEYINPUT57), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n598), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n598), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G164), .B2(G1384), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(G1384), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n983), .B1(new_n896), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1031), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1348), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n896), .A2(new_n974), .A3(new_n1020), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1019), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1025), .B1(new_n1024), .B2(new_n974), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n978), .A2(new_n1019), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(G2067), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n983), .B1(new_n978), .B2(new_n1020), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1348), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1052), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1054), .A2(new_n1059), .A3(new_n633), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1038), .B1(new_n1031), .B2(new_n1044), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1045), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT60), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1050), .A2(KEYINPUT120), .A3(new_n1053), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1057), .B2(new_n1052), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n915), .A3(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT60), .B(new_n633), .C1(new_n1054), .C2(new_n1059), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT45), .B1(new_n1024), .B2(new_n974), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1041), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1019), .B1(new_n899), .B2(new_n1071), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1070), .A2(new_n1072), .A3(G1996), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1051), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n1076), .B2(new_n579), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1078), .B(new_n578), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1069), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1031), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1061), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1031), .A2(new_n1044), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1038), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(KEYINPUT61), .A3(new_n1045), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1062), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n748), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n443), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  OAI21_X1  g668(.A(G2105), .B1(new_n487), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1018), .A2(KEYINPUT122), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n479), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n896), .B2(new_n1041), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n980), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1040), .A2(KEYINPUT114), .A3(new_n1042), .ZN(new_n1101));
  AOI21_X1  g676(.A(G2078), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1091), .B(new_n1098), .C1(new_n1102), .C2(KEYINPUT53), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  AOI21_X1  g679(.A(G301), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n983), .B1(new_n975), .B2(new_n1039), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1024), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1091), .C1(new_n1102), .C2(KEYINPUT53), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1107), .B1(new_n1112), .B2(G301), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(G301), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1103), .A2(G171), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1981), .ZN(new_n1118));
  XNOR2_X1  g693(.A(G305), .B(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT49), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT49), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n812), .A2(new_n1118), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G305), .A2(G1981), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(new_n1124), .A3(G8), .A4(new_n1051), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n608), .A2(G1976), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(G8), .A3(new_n1051), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT52), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n608), .B2(G1976), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1125), .B(new_n1128), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G8), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1100), .A2(new_n809), .A3(new_n1101), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1055), .A2(new_n1056), .A3(new_n796), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(G303), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G166), .A2(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(KEYINPUT55), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT116), .B1(new_n1137), .B2(KEYINPUT55), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1019), .B1(new_n978), .B2(new_n1020), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n796), .A3(new_n1026), .A4(new_n1021), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G8), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1140), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n740), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1055), .A2(new_n1056), .A3(new_n787), .ZN(new_n1152));
  OAI21_X1  g727(.A(G286), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1109), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1019), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n740), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1055), .A2(new_n1056), .A3(new_n787), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(G168), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(G8), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(G8), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(KEYINPUT51), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1132), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT51), .B1(new_n1164), .B2(KEYINPUT121), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1158), .A2(G8), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1149), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1090), .A2(new_n1114), .A3(new_n1117), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G288), .A2(G1976), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1125), .A2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(G8), .B(new_n1051), .C1(new_n1171), .C2(new_n1123), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1132), .B(new_n1140), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1174), .B2(new_n1131), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1142), .A2(new_n1148), .A3(G171), .A4(new_n1111), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1163), .A2(new_n1167), .A3(new_n1176), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1160), .A2(new_n1182), .A3(G286), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1142), .B(new_n1183), .C1(new_n1141), .C2(new_n1135), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1141), .B1(new_n1146), .B2(G8), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1185), .A2(new_n1173), .A3(new_n1131), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1160), .A2(G286), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT118), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1142), .A2(new_n1148), .A3(KEYINPUT118), .A4(new_n1187), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1182), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1184), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1169), .A2(new_n1181), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n1193));
  NAND2_X1  g768(.A1(G290), .A2(G1986), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n985), .B1(new_n987), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1000), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1193), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1012), .B1(new_n1197), .B2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g774(.A1(G227), .A2(new_n465), .ZN(new_n1201));
  NOR3_X1   g775(.A1(G229), .A2(G401), .A3(new_n1201), .ZN(new_n1202));
  AND3_X1   g776(.A1(new_n1202), .A2(new_n970), .A3(new_n910), .ZN(G308));
  NAND3_X1  g777(.A1(new_n1202), .A2(new_n970), .A3(new_n910), .ZN(G225));
endmodule


