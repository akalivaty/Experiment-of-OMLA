

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U557 ( .A1(n715), .A2(n714), .ZN(n756) );
  INV_X2 U558 ( .A(n756), .ZN(n751) );
  INV_X1 U559 ( .A(KEYINPUT95), .ZN(n759) );
  XNOR2_X1 U560 ( .A(n759), .B(KEYINPUT30), .ZN(n760) );
  XNOR2_X1 U561 ( .A(n761), .B(n760), .ZN(n762) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n749) );
  XNOR2_X1 U563 ( .A(n750), .B(n749), .ZN(n755) );
  NAND2_X1 U564 ( .A1(G8), .A2(n756), .ZN(n795) );
  NOR2_X1 U565 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U566 ( .A1(G651), .A2(n628), .ZN(n644) );
  NOR2_X2 U567 ( .A1(n572), .A2(n571), .ZN(n1007) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U569 ( .A1(n641), .A2(G89), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n522), .B(KEYINPUT4), .ZN(n525) );
  INV_X1 U571 ( .A(G651), .ZN(n527) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  OR2_X1 U573 ( .A1(n527), .A2(n628), .ZN(n523) );
  XNOR2_X2 U574 ( .A(KEYINPUT65), .B(n523), .ZN(n640) );
  NAND2_X1 U575 ( .A1(G76), .A2(n640), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U577 ( .A(KEYINPUT5), .B(n526), .ZN(n535) );
  NOR2_X1 U578 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n528), .Z(n529) );
  XNOR2_X1 U580 ( .A(KEYINPUT66), .B(n529), .ZN(n645) );
  NAND2_X1 U581 ( .A1(G63), .A2(n645), .ZN(n530) );
  XOR2_X1 U582 ( .A(KEYINPUT77), .B(n530), .Z(n532) );
  NAND2_X1 U583 ( .A1(n644), .A2(G51), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U587 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  XOR2_X1 U588 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X2 U590 ( .A(KEYINPUT17), .B(n537), .Z(n894) );
  NAND2_X1 U591 ( .A1(n894), .A2(G137), .ZN(n545) );
  INV_X1 U592 ( .A(G2104), .ZN(n540) );
  AND2_X1 U593 ( .A1(n540), .A2(G2105), .ZN(n888) );
  NAND2_X1 U594 ( .A1(G125), .A2(n888), .ZN(n539) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U596 ( .A1(G113), .A2(n886), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n543) );
  NOR2_X4 U598 ( .A1(G2105), .A2(n540), .ZN(n892) );
  NAND2_X1 U599 ( .A1(G101), .A2(n892), .ZN(n541) );
  XNOR2_X1 U600 ( .A(KEYINPUT23), .B(n541), .ZN(n542) );
  NOR2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U603 ( .A(KEYINPUT64), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n547), .B(n546), .ZN(G160) );
  NAND2_X1 U605 ( .A1(n640), .A2(G77), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT68), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G90), .A2(n641), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT9), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G52), .A2(n644), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G64), .A2(n645), .ZN(n554) );
  XNOR2_X1 U613 ( .A(KEYINPUT67), .B(n554), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  NAND2_X1 U617 ( .A1(G94), .A2(G452), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n560) );
  INV_X1 U622 ( .A(G223), .ZN(n820) );
  NAND2_X1 U623 ( .A1(G567), .A2(n820), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(G234) );
  NAND2_X1 U625 ( .A1(n645), .A2(G56), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT73), .B(n561), .Z(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT14), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G43), .A2(n644), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n641), .A2(G81), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n565), .Z(n568) );
  NAND2_X1 U632 ( .A1(n640), .A2(G68), .ZN(n566) );
  XOR2_X1 U633 ( .A(n566), .B(KEYINPUT74), .Z(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT75), .B(n569), .Z(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n1007), .A2(G860), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G79), .A2(n640), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G54), .A2(n644), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G92), .A2(n641), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G66), .A2(n645), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U646 ( .A(KEYINPUT76), .B(n577), .ZN(n578) );
  NOR2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT15), .ZN(n998) );
  INV_X1 U649 ( .A(G868), .ZN(n595) );
  NAND2_X1 U650 ( .A1(n998), .A2(n595), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G78), .A2(n640), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G91), .A2(n641), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n644), .A2(G53), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G65), .A2(n645), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U659 ( .A(KEYINPUT70), .B(n589), .Z(G299) );
  NOR2_X1 U660 ( .A1(G286), .A2(n595), .ZN(n591) );
  NOR2_X1 U661 ( .A1(G299), .A2(G868), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(G297) );
  INV_X1 U663 ( .A(G860), .ZN(n610) );
  NAND2_X1 U664 ( .A1(n610), .A2(G559), .ZN(n592) );
  INV_X1 U665 ( .A(n998), .ZN(n608) );
  NAND2_X1 U666 ( .A1(n592), .A2(n608), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U668 ( .A1(n608), .A2(G868), .ZN(n594) );
  NOR2_X1 U669 ( .A1(G559), .A2(n594), .ZN(n597) );
  AND2_X1 U670 ( .A1(n595), .A2(n1007), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n888), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G99), .A2(n892), .ZN(n599) );
  XNOR2_X1 U675 ( .A(n599), .B(KEYINPUT78), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G135), .A2(n894), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G111), .A2(n886), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n922) );
  XNOR2_X1 U681 ( .A(n922), .B(G2096), .ZN(n607) );
  INV_X1 U682 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(n1007), .ZN(n656) );
  NAND2_X1 U686 ( .A1(n610), .A2(n656), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G67), .A2(n645), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT79), .B(n611), .Z(n613) );
  NAND2_X1 U689 ( .A1(n644), .A2(G55), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U691 ( .A(KEYINPUT80), .B(n614), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G80), .A2(n640), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G93), .A2(n641), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n658) );
  XOR2_X1 U696 ( .A(n619), .B(n658), .Z(G145) );
  NAND2_X1 U697 ( .A1(G73), .A2(n640), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G86), .A2(n641), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G61), .A2(n645), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G48), .A2(n644), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT81), .B(n623), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U706 ( .A1(G87), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n645), .A2(n631), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n644), .A2(G49), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(G288) );
  AND2_X1 U712 ( .A1(n640), .A2(G72), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G85), .A2(n641), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G60), .A2(n645), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n644), .A2(G47), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G75), .A2(n640), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G88), .A2(n641), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n644), .A2(G50), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G62), .A2(n645), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(G166) );
  XNOR2_X1 U726 ( .A(KEYINPUT19), .B(G305), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n650), .B(G288), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n658), .B(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(G290), .B(G166), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U731 ( .A(G299), .ZN(n744) );
  XNOR2_X1 U732 ( .A(n654), .B(n744), .ZN(n907) );
  XOR2_X1 U733 ( .A(n907), .B(KEYINPUT82), .Z(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(G868), .ZN(n660) );
  OR2_X1 U736 ( .A1(G868), .A2(n658), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n662), .ZN(n664) );
  XOR2_X1 U741 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n663) );
  XNOR2_X1 U742 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U743 ( .A1(G2072), .A2(n665), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U745 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U746 ( .A1(G219), .A2(G220), .ZN(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NOR2_X1 U750 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G96), .A2(n670), .ZN(n826) );
  NAND2_X1 U752 ( .A1(n826), .A2(G2106), .ZN(n674) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U754 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U755 ( .A1(G108), .A2(n672), .ZN(n827) );
  NAND2_X1 U756 ( .A1(n827), .A2(G567), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n674), .A2(n673), .ZN(n828) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U759 ( .A1(n828), .A2(n675), .ZN(n825) );
  NAND2_X1 U760 ( .A1(n825), .A2(G36), .ZN(n676) );
  XNOR2_X1 U761 ( .A(KEYINPUT86), .B(n676), .ZN(G176) );
  NAND2_X1 U762 ( .A1(G102), .A2(n892), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G138), .A2(n894), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G126), .A2(n888), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G114), .A2(n886), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U770 ( .A(G1986), .B(G290), .ZN(n1018) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n684) );
  XNOR2_X1 U773 ( .A(KEYINPUT87), .B(n684), .ZN(n714) );
  INV_X1 U774 ( .A(n714), .ZN(n685) );
  NOR2_X1 U775 ( .A1(n715), .A2(n685), .ZN(n815) );
  NAND2_X1 U776 ( .A1(n1018), .A2(n815), .ZN(n804) );
  NAND2_X1 U777 ( .A1(G119), .A2(n888), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G107), .A2(n886), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U780 ( .A1(G95), .A2(n892), .ZN(n688) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(n688), .ZN(n689) );
  NOR2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n894), .A2(G131), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n870) );
  NAND2_X1 U785 ( .A1(G1991), .A2(n870), .ZN(n701) );
  NAND2_X1 U786 ( .A1(G129), .A2(n888), .ZN(n694) );
  NAND2_X1 U787 ( .A1(G117), .A2(n886), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n892), .A2(G105), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n695), .Z(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n894), .A2(G141), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n873) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n873), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n925) );
  NAND2_X1 U796 ( .A1(n925), .A2(n815), .ZN(n702) );
  XOR2_X1 U797 ( .A(KEYINPUT90), .B(n702), .Z(n807) );
  INV_X1 U798 ( .A(n807), .ZN(n713) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n703) );
  XNOR2_X1 U800 ( .A(n703), .B(KEYINPUT88), .ZN(n813) );
  NAND2_X1 U801 ( .A1(G104), .A2(n892), .ZN(n705) );
  NAND2_X1 U802 ( .A1(G140), .A2(n894), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U804 ( .A(KEYINPUT34), .B(n706), .ZN(n711) );
  NAND2_X1 U805 ( .A1(G128), .A2(n888), .ZN(n708) );
  NAND2_X1 U806 ( .A1(G116), .A2(n886), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U808 ( .A(KEYINPUT35), .B(n709), .Z(n710) );
  NOR2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U810 ( .A(KEYINPUT36), .B(n712), .ZN(n902) );
  NOR2_X1 U811 ( .A1(n813), .A2(n902), .ZN(n929) );
  NAND2_X1 U812 ( .A1(n815), .A2(n929), .ZN(n811) );
  NAND2_X1 U813 ( .A1(n713), .A2(n811), .ZN(n802) );
  NOR2_X1 U814 ( .A1(G1981), .A2(G305), .ZN(n716) );
  XOR2_X1 U815 ( .A(n716), .B(KEYINPUT24), .Z(n717) );
  NOR2_X1 U816 ( .A1(n795), .A2(n717), .ZN(n800) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NAND2_X1 U818 ( .A1(n785), .A2(KEYINPUT33), .ZN(n718) );
  NOR2_X1 U819 ( .A1(n795), .A2(n718), .ZN(n790) );
  XNOR2_X1 U820 ( .A(KEYINPUT93), .B(G1341), .ZN(n720) );
  INV_X1 U821 ( .A(KEYINPUT26), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n751), .A2(n726), .ZN(n719) );
  NAND2_X1 U823 ( .A1(n720), .A2(n719), .ZN(n725) );
  INV_X1 U824 ( .A(KEYINPUT93), .ZN(n723) );
  INV_X1 U825 ( .A(G1996), .ZN(n956) );
  NOR2_X1 U826 ( .A1(n956), .A2(n726), .ZN(n721) );
  NOR2_X1 U827 ( .A1(n756), .A2(n721), .ZN(n722) );
  NAND2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U830 ( .A1(n956), .A2(n726), .ZN(n727) );
  NAND2_X1 U831 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U832 ( .A(KEYINPUT94), .B(n729), .ZN(n734) );
  NAND2_X1 U833 ( .A1(G1348), .A2(n756), .ZN(n731) );
  NAND2_X1 U834 ( .A1(G2067), .A2(n751), .ZN(n730) );
  NAND2_X1 U835 ( .A1(n731), .A2(n730), .ZN(n735) );
  NAND2_X1 U836 ( .A1(n998), .A2(n735), .ZN(n732) );
  NAND2_X1 U837 ( .A1(n1007), .A2(n732), .ZN(n733) );
  NOR2_X1 U838 ( .A1(n734), .A2(n733), .ZN(n737) );
  NOR2_X1 U839 ( .A1(n735), .A2(n998), .ZN(n736) );
  NOR2_X1 U840 ( .A1(n737), .A2(n736), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n751), .A2(G2072), .ZN(n738) );
  XNOR2_X1 U842 ( .A(KEYINPUT27), .B(n738), .ZN(n741) );
  XOR2_X1 U843 ( .A(KEYINPUT91), .B(G1956), .Z(n983) );
  NAND2_X1 U844 ( .A1(n983), .A2(n756), .ZN(n739) );
  XOR2_X1 U845 ( .A(KEYINPUT92), .B(n739), .Z(n740) );
  NOR2_X1 U846 ( .A1(n741), .A2(n740), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n745), .A2(n744), .ZN(n742) );
  NAND2_X1 U848 ( .A1(n743), .A2(n742), .ZN(n748) );
  NOR2_X1 U849 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U850 ( .A(n746), .B(KEYINPUT28), .Z(n747) );
  NAND2_X1 U851 ( .A1(n748), .A2(n747), .ZN(n750) );
  OR2_X1 U852 ( .A1(n751), .A2(G1961), .ZN(n753) );
  XNOR2_X1 U853 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U854 ( .A1(n751), .A2(n955), .ZN(n752) );
  NAND2_X1 U855 ( .A1(n753), .A2(n752), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n763), .A2(G171), .ZN(n754) );
  NAND2_X1 U857 ( .A1(n755), .A2(n754), .ZN(n768) );
  NOR2_X1 U858 ( .A1(G1966), .A2(n795), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G2084), .A2(n756), .ZN(n776) );
  INV_X1 U860 ( .A(n776), .ZN(n757) );
  NAND2_X1 U861 ( .A1(G8), .A2(n757), .ZN(n758) );
  OR2_X1 U862 ( .A1(n777), .A2(n758), .ZN(n761) );
  NOR2_X1 U863 ( .A1(G168), .A2(n762), .ZN(n765) );
  NOR2_X1 U864 ( .A1(G171), .A2(n763), .ZN(n764) );
  NOR2_X1 U865 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U866 ( .A(KEYINPUT31), .B(n766), .Z(n767) );
  NAND2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n778), .A2(G286), .ZN(n773) );
  NOR2_X1 U869 ( .A1(G1971), .A2(n795), .ZN(n770) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n756), .ZN(n769) );
  NOR2_X1 U871 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U872 ( .A1(n771), .A2(G303), .ZN(n772) );
  NAND2_X1 U873 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U874 ( .A1(n774), .A2(G8), .ZN(n775) );
  XNOR2_X1 U875 ( .A(n775), .B(KEYINPUT32), .ZN(n783) );
  NAND2_X1 U876 ( .A1(G8), .A2(n776), .ZN(n781) );
  INV_X1 U877 ( .A(n778), .ZN(n779) );
  NOR2_X1 U878 ( .A1(n777), .A2(n779), .ZN(n780) );
  NAND2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n794) );
  NOR2_X1 U881 ( .A1(G1971), .A2(G303), .ZN(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n1016) );
  NAND2_X1 U883 ( .A1(n794), .A2(n1016), .ZN(n786) );
  NAND2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  NAND2_X1 U885 ( .A1(n786), .A2(n1012), .ZN(n787) );
  NOR2_X1 U886 ( .A1(n795), .A2(n787), .ZN(n788) );
  NOR2_X1 U887 ( .A1(KEYINPUT33), .A2(n788), .ZN(n789) );
  NOR2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U889 ( .A(G1981), .B(G305), .Z(n1002) );
  NAND2_X1 U890 ( .A1(n791), .A2(n1002), .ZN(n798) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U892 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n818) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n870), .ZN(n923) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n923), .A2(n805), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n873), .ZN(n920) );
  NOR2_X1 U903 ( .A1(n808), .A2(n920), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(KEYINPUT96), .ZN(n810) );
  XNOR2_X1 U905 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n813), .A2(n902), .ZN(n937) );
  NAND2_X1 U908 ( .A1(n814), .A2(n937), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U911 ( .A(n819), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n820), .ZN(G217) );
  INV_X1 U913 ( .A(G661), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G2), .A2(G15), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT98), .B(n823), .Z(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U919 ( .A(G96), .B(KEYINPUT99), .ZN(G221) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  INV_X1 U925 ( .A(n828), .ZN(G319) );
  XNOR2_X1 U926 ( .A(G1341), .B(G2454), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n829), .B(G2430), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(G1348), .ZN(n836) );
  XOR2_X1 U929 ( .A(G2443), .B(G2427), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2438), .B(G2446), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n834) );
  XOR2_X1 U932 ( .A(G2451), .B(G2435), .Z(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n837), .A2(G14), .ZN(n838) );
  XNOR2_X1 U936 ( .A(KEYINPUT97), .B(n838), .ZN(G401) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2678), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2096), .B(G2100), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U946 ( .A(G2078), .B(G2084), .Z(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1956), .B(G1961), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n860) );
  XOR2_X1 U951 ( .A(KEYINPUT104), .B(G2474), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1976), .B(KEYINPUT102), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(G1981), .B(G1971), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT103), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n888), .A2(G124), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G136), .A2(n894), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT105), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G112), .A2(n886), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n892), .A2(G100), .ZN(n867) );
  XOR2_X1 U969 ( .A(KEYINPUT106), .B(n867), .Z(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(G162) );
  XNOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n870), .B(KEYINPUT110), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n922), .B(G160), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n876), .B(n875), .Z(n878) );
  XNOR2_X1 U977 ( .A(G164), .B(G162), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n904) );
  NAND2_X1 U979 ( .A1(G130), .A2(n888), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n886), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G106), .A2(n892), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G142), .A2(n894), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n900) );
  NAND2_X1 U987 ( .A1(n886), .A2(G115), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT109), .B(n887), .Z(n890) );
  NAND2_X1 U989 ( .A1(n888), .A2(G127), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .ZN(n899) );
  NAND2_X1 U992 ( .A1(n892), .A2(G103), .ZN(n893) );
  XOR2_X1 U993 ( .A(KEYINPUT107), .B(n893), .Z(n896) );
  NAND2_X1 U994 ( .A1(n894), .A2(G139), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(KEYINPUT108), .B(n897), .Z(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n932) );
  XNOR2_X1 U998 ( .A(n900), .B(n932), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(n906) );
  XOR2_X1 U1002 ( .A(KEYINPUT111), .B(n906), .Z(G395) );
  XNOR2_X1 U1003 ( .A(n907), .B(KEYINPUT112), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n998), .B(G286), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1006 ( .A(n1007), .B(G171), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(KEYINPUT49), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n914), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT113), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n921), .Z(n931) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n940) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n935) );
  XNOR2_X1 U1028 ( .A(KEYINPUT114), .B(n932), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n933), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(n936), .B(KEYINPUT50), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1038 ( .A(G29), .B(KEYINPUT119), .ZN(n968) );
  XOR2_X1 U1039 ( .A(G2090), .B(G35), .Z(n948) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT118), .B(n945), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(n946), .B(KEYINPUT54), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n965) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1045 ( .A1(G28), .A2(n949), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n950), .B(KEYINPUT115), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n961) );
  XOR2_X1 U1051 ( .A(n955), .B(G27), .Z(n958) );
  XOR2_X1 U1052 ( .A(n956), .B(G32), .Z(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1054 ( .A(n959), .B(KEYINPUT116), .Z(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT53), .B(n962), .Z(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT117), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n969), .ZN(n1026) );
  XOR2_X1 U1062 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n977) );
  XNOR2_X1 U1063 ( .A(G1986), .B(G24), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G1976), .B(G23), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(KEYINPUT58), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n977), .B(n976), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G5), .B(G1961), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n992) );
  XOR2_X1 U1075 ( .A(G1348), .B(KEYINPUT59), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G4), .B(n982), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G20), .B(n983), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G1981), .B(G6), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(n993), .B(KEYINPUT61), .Z(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G16), .B(KEYINPUT122), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(n997), .ZN(n1024) );
  XNOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .ZN(n1022) );
  XNOR2_X1 U1091 ( .A(G301), .B(G1961), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n998), .B(G1348), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1001), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(n1004), .B(KEYINPUT57), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1341), .B(n1007), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(KEYINPUT121), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1020) );
  NAND2_X1 U1102 ( .A1(G1971), .A2(G303), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(G1956), .B(G299), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

