//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n441, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(G124), .A2(new_n474), .B1(new_n465), .B2(G136), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n475), .A2(new_n479), .ZN(G162));
  OAI21_X1  g055(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(G114), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT70), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT69), .A2(G114), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT69), .A2(G114), .ZN(new_n486));
  OAI211_X1 g061(.A(KEYINPUT70), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n482), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n473), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G138), .A4(new_n473), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n492), .A2(G126), .A3(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n510), .A2(new_n517), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n507), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n510), .A2(new_n529), .B1(new_n512), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n507), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT71), .B(G81), .Z(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n510), .A2(new_n535), .B1(new_n512), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT72), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G188));
  NAND3_X1  g120(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT9), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G91), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n507), .B1(new_n510), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT73), .ZN(G299));
  INV_X1    g128(.A(G171), .ZN(G301));
  INV_X1    g129(.A(G168), .ZN(G286));
  OAI21_X1  g130(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n505), .A2(new_n509), .A3(G87), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  INV_X1    g134(.A(new_n512), .ZN(new_n560));
  NAND2_X1  g135(.A1(G73), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n504), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(G48), .A2(new_n560), .B1(new_n563), .B2(G651), .ZN(new_n564));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(new_n510), .ZN(G305));
  INV_X1    g141(.A(G85), .ZN(new_n567));
  INV_X1    g142(.A(G47), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n510), .A2(new_n567), .B1(new_n512), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n507), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G171), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G92), .ZN(new_n579));
  OR3_X1    g154(.A1(new_n510), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n510), .B2(new_n579), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n560), .A2(G54), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n507), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT10), .B1(new_n580), .B2(new_n581), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n578), .B1(new_n587), .B2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(KEYINPUT75), .B2(new_n577), .ZN(G321));
  XOR2_X1   g165(.A(G321), .B(KEYINPUT77), .Z(G284));
  NAND2_X1  g166(.A1(G299), .A2(new_n576), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n576), .B2(G168), .ZN(G297));
  OAI21_X1  g168(.A(new_n592), .B1(new_n576), .B2(G168), .ZN(G280));
  XOR2_X1   g169(.A(KEYINPUT78), .B(G559), .Z(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n587), .B1(G860), .B2(new_n596), .ZN(G148));
  OAI21_X1  g172(.A(new_n576), .B1(new_n534), .B2(new_n537), .ZN(new_n598));
  INV_X1    g173(.A(new_n587), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n595), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n600), .B2(new_n576), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n492), .A2(new_n466), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT13), .Z(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(G2100), .ZN(new_n606));
  AOI22_X1  g181(.A1(G123), .A2(new_n474), .B1(new_n465), .B2(G135), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n473), .A2(KEYINPUT79), .A3(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n473), .B2(G111), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n605), .A2(G2100), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n606), .A2(new_n612), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(KEYINPUT15), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2435), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2427), .B(G2438), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G1341), .B(G1348), .Z(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT81), .ZN(new_n630));
  OAI21_X1  g205(.A(G14), .B1(new_n626), .B2(new_n628), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(new_n631), .ZN(G401));
  XOR2_X1   g207(.A(G2072), .B(G2078), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT17), .ZN(new_n634));
  XOR2_X1   g209(.A(G2067), .B(G2678), .Z(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n635), .B2(new_n633), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n636), .B1(KEYINPUT82), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(KEYINPUT82), .B2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n637), .A3(new_n635), .ZN(new_n641));
  INV_X1    g216(.A(new_n637), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n642), .A2(new_n635), .A3(new_n633), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n640), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(G2096), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n652), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT84), .ZN(new_n656));
  OR3_X1    g231(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT84), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n659));
  OAI221_X1 g234(.A(new_n653), .B1(new_n650), .B2(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n658), .B2(new_n659), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G1991), .ZN(new_n662));
  INV_X1    g237(.A(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G1986), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT86), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G22), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(G166), .B2(new_n671), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(G1971), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(G6), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G305), .B2(G16), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT32), .B(G1981), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(G1971), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n674), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR2_X1   g256(.A1(G16), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g258(.A1(G288), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n556), .A2(new_n558), .A3(new_n557), .A4(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n686), .B2(G16), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n680), .A2(new_n681), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT34), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n671), .A2(G24), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n574), .B2(new_n671), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n474), .A2(G119), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n465), .A2(G131), .ZN(new_n699));
  OR2_X1    g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n697), .B1(new_n703), .B2(new_n696), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n691), .A2(new_n695), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT36), .Z(new_n708));
  INV_X1    g283(.A(KEYINPUT23), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n671), .A2(G20), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n709), .B(new_n710), .C1(G299), .C2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1956), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n671), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n671), .ZN(new_n716));
  INV_X1    g291(.A(G1966), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G5), .A2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G171), .B2(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G1961), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n611), .A2(new_n696), .ZN(new_n722));
  INV_X1    g297(.A(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n718), .A2(new_n721), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NOR2_X1   g305(.A1(G164), .A2(new_n696), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G27), .B2(new_n696), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n696), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n696), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT29), .Z(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n734), .B(new_n740), .C1(new_n739), .C2(new_n738), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n473), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n466), .A2(G103), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT92), .Z(new_n746));
  AOI22_X1  g321(.A1(new_n746), .A2(KEYINPUT25), .B1(G139), .B2(new_n465), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n747), .C1(KEYINPUT25), .C2(new_n746), .ZN(new_n748));
  MUX2_X1   g323(.A(G33), .B(new_n748), .S(G29), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2072), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G32), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n474), .A2(G129), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n466), .A2(G105), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(G141), .C2(new_n465), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G34), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G160), .B2(G29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G2084), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G2084), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G1961), .B2(new_n720), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n750), .A2(new_n762), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n714), .A2(new_n730), .A3(new_n741), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n671), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n587), .B2(new_n671), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT89), .B(G1348), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n696), .A2(G26), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n465), .A2(G140), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n474), .A2(G128), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n779), .A2(G104), .A3(G2105), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(G104), .B2(G2105), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n473), .A2(G116), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n780), .A2(new_n781), .A3(G2104), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n777), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n776), .B1(new_n785), .B2(new_n696), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n776), .B(new_n786), .S(KEYINPUT28), .Z(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G2067), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n671), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n538), .B2(new_n671), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n775), .A2(new_n788), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n708), .A2(new_n771), .A3(new_n794), .ZN(G311));
  INV_X1    g370(.A(G311), .ZN(G150));
  NAND2_X1  g371(.A1(new_n587), .A2(G559), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n507), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  INV_X1    g377(.A(G55), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n510), .A2(new_n802), .B1(new_n512), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n538), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n799), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n805), .A2(new_n809), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT97), .Z(G145));
  XNOR2_X1  g390(.A(new_n785), .B(new_n498), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n748), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n759), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n465), .A2(G142), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n473), .A2(G118), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n474), .A2(G130), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n702), .B(new_n604), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT99), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(KEYINPUT99), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n818), .A2(new_n828), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n611), .B(G160), .Z(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G162), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND4_X1   g410(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n832), .B2(new_n829), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n836), .A2(G37), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(G395));
  XOR2_X1   g415(.A(new_n574), .B(new_n686), .Z(new_n841));
  XNOR2_X1  g416(.A(G303), .B(G305), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT42), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n600), .B(new_n807), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n599), .B(G299), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(KEYINPUT41), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n845), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n844), .B(new_n849), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G868), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G868), .B2(new_n805), .ZN(G331));
  XOR2_X1   g427(.A(G331), .B(KEYINPUT101), .Z(G295));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n854));
  XNOR2_X1  g429(.A(G171), .B(G168), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n806), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n846), .A2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n854), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n843), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n864), .B2(new_n843), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT43), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n843), .B1(new_n859), .B2(new_n860), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n871));
  OAI211_X1 g446(.A(new_n867), .B(KEYINPUT44), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n873), .A3(new_n871), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n866), .B2(new_n871), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(G397));
  INV_X1    g454(.A(G1384), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n498), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT45), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(G160), .A2(G40), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n663), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT124), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT46), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(KEYINPUT46), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G2067), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n784), .B(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n759), .B(new_n892), .C1(G1996), .C2(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n885), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT125), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT47), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n892), .B1(new_n759), .B2(new_n663), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n758), .A2(G1996), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT106), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n702), .B(new_n705), .Z(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n885), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(G290), .A2(G1986), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n885), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT48), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n703), .A2(new_n705), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n901), .A2(new_n907), .B1(G2067), .B2(new_n784), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n903), .A2(new_n906), .B1(new_n908), .B2(new_n885), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT123), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT115), .ZN(new_n912));
  INV_X1    g487(.A(G8), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n880), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n884), .B1(new_n914), .B2(KEYINPUT108), .ZN(new_n915));
  OAI21_X1  g490(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT70), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n487), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n496), .B1(new_n919), .B2(new_n482), .ZN(new_n920));
  AOI21_X1  g495(.A(G1384), .B1(new_n920), .B2(new_n495), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT45), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n921), .B2(KEYINPUT45), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n881), .A2(new_n925), .A3(new_n882), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(new_n923), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1971), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  AOI211_X1 g505(.A(KEYINPUT109), .B(G1384), .C1(new_n920), .C2(new_n495), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n498), .B2(new_n880), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n884), .B1(KEYINPUT50), .B2(new_n881), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n739), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n913), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g512(.A1(G303), .A2(G8), .B1(KEYINPUT110), .B2(KEYINPUT55), .ZN(new_n938));
  OR2_X1    g513(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n938), .B(new_n939), .Z(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n931), .A2(new_n933), .A3(KEYINPUT45), .ZN(new_n942));
  INV_X1    g517(.A(new_n884), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n914), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n717), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G2084), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n934), .A2(new_n946), .A3(new_n935), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n881), .A2(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n921), .A2(new_n932), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n884), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n913), .ZN(new_n954));
  INV_X1    g529(.A(G1976), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n684), .B2(new_n685), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT52), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n955), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1981), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(G86), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n505), .A2(new_n509), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n564), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT113), .B1(G305), .B2(G1981), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(KEYINPUT114), .B2(KEYINPUT49), .ZN(new_n970));
  NOR2_X1   g545(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n971), .B(new_n967), .C1(new_n968), .C2(new_n965), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n954), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n959), .A2(new_n961), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n937), .A2(new_n940), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n912), .B1(new_n950), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n940), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n931), .A2(new_n933), .A3(new_n930), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n943), .B1(new_n881), .B2(KEYINPUT50), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(new_n980), .A3(G2090), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n928), .B2(new_n927), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n982), .B2(new_n913), .ZN(new_n983));
  INV_X1    g558(.A(new_n947), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n951), .A2(new_n952), .A3(new_n882), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n884), .B1(KEYINPUT45), .B2(new_n921), .ZN(new_n986));
  AOI21_X1  g561(.A(G1966), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(G8), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G286), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n974), .A2(new_n983), .A3(new_n975), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n959), .A2(new_n973), .A3(new_n961), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n940), .B2(new_n937), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n941), .A2(new_n949), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(KEYINPUT115), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n977), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G288), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n973), .A2(new_n955), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(G305), .A2(G1981), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n975), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1002), .A2(new_n954), .B1(new_n1003), .B2(new_n974), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n913), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n988), .A2(KEYINPUT51), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1009), .B(G8), .C1(new_n948), .C2(G286), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n948), .A2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1008), .A2(new_n1010), .A3(new_n1014), .A4(new_n1011), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT121), .B(G1961), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n934), .B2(new_n935), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n925), .B1(new_n881), .B2(new_n882), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT107), .B(KEYINPUT45), .C1(new_n498), .C2(new_n880), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(new_n733), .A3(new_n923), .A4(new_n915), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(G2078), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n985), .A2(new_n986), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G301), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1013), .A2(new_n1015), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n927), .B2(G2078), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1018), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1032), .A2(new_n923), .A3(new_n943), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n883), .A3(new_n1025), .ZN(new_n1034));
  AND4_X1   g609(.A1(G301), .A2(new_n1030), .A3(new_n1031), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1029), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1012), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1021), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n713), .B1(new_n979), .B2(new_n980), .ZN(new_n1040));
  NAND2_X1  g615(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1041), .B(new_n1044), .C1(new_n548), .C2(new_n551), .ZN(new_n1045));
  INV_X1    g620(.A(new_n551), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n1042), .A3(new_n1043), .A4(new_n547), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(new_n1040), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(KEYINPUT117), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n934), .A2(new_n935), .ZN(new_n1056));
  INV_X1    g631(.A(G1348), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1057), .B1(new_n891), .B2(new_n953), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1055), .A2(KEYINPUT118), .B1(new_n599), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1060), .B(new_n1054), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1050), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT59), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT119), .B(G1996), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT58), .B(G1341), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n927), .A2(new_n1066), .B1(new_n953), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1068), .B2(new_n538), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n538), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n934), .B2(new_n935), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n943), .B(new_n891), .C1(new_n931), .C2(new_n933), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n599), .B1(new_n1058), .B2(KEYINPUT60), .ZN(new_n1079));
  NOR4_X1   g654(.A1(new_n1075), .A2(new_n1077), .A3(new_n1074), .A4(new_n587), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1049), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1050), .B1(new_n1082), .B2(KEYINPUT61), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1039), .A2(new_n1084), .A3(new_n1040), .A4(new_n1049), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1073), .A2(new_n1081), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1037), .B1(new_n1062), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1030), .A2(G301), .A3(new_n1031), .A4(new_n1026), .ZN(new_n1091));
  AND4_X1   g666(.A1(new_n1088), .A2(new_n1090), .A3(KEYINPUT54), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1029), .B1(new_n1089), .B2(G171), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1093), .B2(new_n1091), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1028), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n994), .A2(new_n983), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1005), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(G290), .A2(G1986), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n885), .B1(new_n1099), .B2(new_n904), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n903), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n911), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1069), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1068), .A2(new_n538), .A3(new_n1072), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1083), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1062), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1012), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1024), .A2(G301), .A3(new_n1034), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT54), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1095), .A2(new_n1107), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1013), .A2(new_n1015), .A3(new_n1027), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1097), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n997), .A2(new_n1004), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n911), .B(new_n1101), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n910), .B1(new_n1102), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT126), .B(new_n910), .C1(new_n1102), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g699(.A(G319), .ZN(new_n1126));
  NOR3_X1   g700(.A1(G401), .A2(new_n1126), .A3(G227), .ZN(new_n1127));
  OAI21_X1  g701(.A(new_n669), .B1(new_n1127), .B2(KEYINPUT127), .ZN(new_n1128));
  AND2_X1   g702(.A1(new_n1127), .A2(KEYINPUT127), .ZN(new_n1129));
  NOR3_X1   g703(.A1(new_n1128), .A2(new_n838), .A3(new_n1129), .ZN(new_n1130));
  OAI211_X1 g704(.A(new_n1130), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(G225));
  INV_X1    g705(.A(G225), .ZN(G308));
endmodule


