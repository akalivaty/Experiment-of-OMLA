

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X2 U322 ( .A(n440), .B(n439), .Z(n449) );
  NOR2_X1 U323 ( .A1(n459), .A2(n458), .ZN(n460) );
  BUF_X1 U324 ( .A(n447), .Z(n448) );
  XNOR2_X1 U325 ( .A(n421), .B(n290), .ZN(n337) );
  AND2_X1 U326 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  INV_X1 U327 ( .A(KEYINPUT25), .ZN(n382) );
  XNOR2_X1 U328 ( .A(n382), .B(KEYINPUT94), .ZN(n383) );
  XNOR2_X1 U329 ( .A(n384), .B(n383), .ZN(n388) );
  INV_X1 U330 ( .A(KEYINPUT118), .ZN(n464) );
  XNOR2_X1 U331 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  XNOR2_X1 U332 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U333 ( .A(KEYINPUT48), .B(n460), .Z(n543) );
  XNOR2_X1 U334 ( .A(n468), .B(KEYINPUT119), .ZN(n563) );
  XNOR2_X1 U335 ( .A(n338), .B(n337), .ZN(n346) );
  INV_X1 U336 ( .A(G50GAT), .ZN(n444) );
  XNOR2_X1 U337 ( .A(n470), .B(KEYINPUT122), .ZN(n471) );
  XNOR2_X1 U338 ( .A(n444), .B(KEYINPUT102), .ZN(n445) );
  XNOR2_X1 U339 ( .A(n472), .B(n471), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n446), .B(n445), .ZN(G1331GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n292) );
  XNOR2_X1 U342 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U344 ( .A(n293), .B(KEYINPUT22), .Z(n295) );
  XOR2_X1 U345 ( .A(G141GAT), .B(G22GAT), .Z(n434) );
  XNOR2_X1 U346 ( .A(G50GAT), .B(n434), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n301) );
  XOR2_X1 U348 ( .A(G78GAT), .B(G148GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(G204GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n415) );
  XOR2_X1 U351 ( .A(G211GAT), .B(n415), .Z(n299) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n301), .B(n300), .Z(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT2), .B(G162GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(KEYINPUT3), .B(n304), .Z(n363) );
  XOR2_X1 U359 ( .A(KEYINPUT21), .B(G218GAT), .Z(n306) );
  XNOR2_X1 U360 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U362 ( .A(G197GAT), .B(n307), .Z(n375) );
  XNOR2_X1 U363 ( .A(n363), .B(n375), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n463) );
  XNOR2_X1 U365 ( .A(n463), .B(KEYINPUT28), .ZN(n505) );
  INV_X1 U366 ( .A(n505), .ZN(n520) );
  XOR2_X1 U367 ( .A(G190GAT), .B(G134GAT), .Z(n332) );
  XOR2_X1 U368 ( .A(G85GAT), .B(G92GAT), .Z(n416) );
  XNOR2_X1 U369 ( .A(n332), .B(n416), .ZN(n311) );
  XOR2_X1 U370 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n312), .B(KEYINPUT73), .Z(n317) );
  XOR2_X1 U373 ( .A(G106GAT), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G99GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U376 ( .A(G218GAT), .B(n315), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n319) );
  NAND2_X1 U379 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n328) );
  XOR2_X1 U382 ( .A(G29GAT), .B(KEYINPUT65), .Z(n323) );
  XNOR2_X1 U383 ( .A(G50GAT), .B(G36GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n439) );
  INV_X1 U387 ( .A(n439), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n326), .B(KEYINPUT11), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n447) );
  XOR2_X1 U390 ( .A(n447), .B(KEYINPUT36), .Z(n583) );
  XOR2_X1 U391 ( .A(KEYINPUT81), .B(KEYINPUT78), .Z(n330) );
  XNOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT82), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT20), .Z(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U396 ( .A(KEYINPUT0), .B(G127GAT), .Z(n349) );
  XNOR2_X1 U397 ( .A(n333), .B(n349), .ZN(n334) );
  XOR2_X1 U398 ( .A(n335), .B(n334), .Z(n338) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G71GAT), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n336), .B(G120GAT), .ZN(n421) );
  XOR2_X1 U401 ( .A(G15GAT), .B(G113GAT), .Z(n340) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G43GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n430) );
  XNOR2_X1 U404 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n341), .B(G176GAT), .ZN(n342) );
  XOR2_X1 U406 ( .A(n342), .B(KEYINPUT19), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n379) );
  XNOR2_X1 U409 ( .A(n430), .B(n379), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n502) );
  XNOR2_X1 U411 ( .A(KEYINPUT83), .B(n502), .ZN(n380) );
  XOR2_X1 U412 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n348) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U415 ( .A(G85GAT), .B(KEYINPUT90), .Z(n351) );
  XNOR2_X1 U416 ( .A(G134GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U418 ( .A(n353), .B(n352), .Z(n355) );
  NAND2_X1 U419 ( .A1(G225GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U421 ( .A(G120GAT), .B(G113GAT), .Z(n357) );
  XNOR2_X1 U422 ( .A(G29GAT), .B(G141GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U425 ( .A(KEYINPUT1), .B(G57GAT), .Z(n361) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G148GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n512) );
  XOR2_X1 U430 ( .A(KEYINPUT92), .B(G92GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(G190GAT), .B(G204GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U433 ( .A(G8GAT), .B(G211GAT), .Z(n398) );
  XOR2_X1 U434 ( .A(n368), .B(n398), .Z(n370) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G36GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U437 ( .A(KEYINPUT91), .B(G64GAT), .Z(n372) );
  NAND2_X1 U438 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U440 ( .A(n374), .B(n373), .Z(n377) );
  XNOR2_X1 U441 ( .A(n375), .B(KEYINPUT93), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n514) );
  XNOR2_X1 U444 ( .A(KEYINPUT27), .B(n514), .ZN(n386) );
  OR2_X1 U445 ( .A1(n512), .A2(n386), .ZN(n542) );
  NOR2_X1 U446 ( .A1(n542), .A2(n505), .ZN(n524) );
  NAND2_X1 U447 ( .A1(n380), .A2(n524), .ZN(n392) );
  INV_X1 U448 ( .A(n502), .ZN(n526) );
  NOR2_X1 U449 ( .A1(n526), .A2(n514), .ZN(n381) );
  NOR2_X1 U450 ( .A1(n463), .A2(n381), .ZN(n384) );
  NAND2_X1 U451 ( .A1(n463), .A2(n526), .ZN(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT26), .B(n385), .ZN(n568) );
  NOR2_X1 U453 ( .A1(n386), .A2(n568), .ZN(n387) );
  NOR2_X1 U454 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n389), .B(KEYINPUT95), .ZN(n390) );
  NAND2_X1 U456 ( .A1(n390), .A2(n512), .ZN(n391) );
  NAND2_X1 U457 ( .A1(n392), .A2(n391), .ZN(n393) );
  XOR2_X1 U458 ( .A(KEYINPUT96), .B(n393), .Z(n475) );
  NOR2_X1 U459 ( .A1(n583), .A2(n475), .ZN(n412) );
  XOR2_X1 U460 ( .A(G155GAT), .B(G71GAT), .Z(n395) );
  XNOR2_X1 U461 ( .A(G22GAT), .B(G15GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n411) );
  XOR2_X1 U463 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n397) );
  XNOR2_X1 U464 ( .A(G57GAT), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n414) );
  XOR2_X1 U466 ( .A(n414), .B(n398), .Z(n400) );
  XNOR2_X1 U467 ( .A(G183GAT), .B(G127GAT), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U469 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n402) );
  NAND2_X1 U470 ( .A1(G231GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U472 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U473 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n406) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G78GAT), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT12), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n551) );
  NAND2_X1 U479 ( .A1(n412), .A2(n551), .ZN(n413) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(n413), .ZN(n511) );
  XOR2_X1 U481 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n425) );
  XOR2_X1 U483 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n423) );
  XOR2_X1 U484 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n419) );
  XNOR2_X1 U485 ( .A(G176GAT), .B(KEYINPUT69), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n427) );
  NAND2_X1 U490 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n574) );
  XOR2_X1 U492 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n429) );
  XNOR2_X1 U493 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n430), .B(G1GAT), .ZN(n432) );
  AND2_X1 U496 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n433), .B(G8GAT), .ZN(n436) );
  XOR2_X1 U499 ( .A(G197GAT), .B(n434), .Z(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n440) );
  INV_X1 U502 ( .A(n449), .ZN(n541) );
  XNOR2_X1 U503 ( .A(KEYINPUT67), .B(n541), .ZN(n555) );
  NAND2_X1 U504 ( .A1(n574), .A2(n555), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n441), .B(KEYINPUT71), .ZN(n477) );
  NAND2_X1 U506 ( .A1(n511), .A2(n477), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n442), .B(KEYINPUT38), .ZN(n443) );
  XNOR2_X1 U508 ( .A(KEYINPUT100), .B(n443), .ZN(n490) );
  NOR2_X1 U509 ( .A1(n520), .A2(n490), .ZN(n446) );
  INV_X1 U510 ( .A(n514), .ZN(n500) );
  XNOR2_X1 U511 ( .A(KEYINPUT41), .B(n574), .ZN(n558) );
  NAND2_X1 U512 ( .A1(n449), .A2(n558), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n450), .B(KEYINPUT46), .ZN(n451) );
  XNOR2_X1 U514 ( .A(KEYINPUT110), .B(n551), .ZN(n535) );
  NAND2_X1 U515 ( .A1(n451), .A2(n535), .ZN(n452) );
  NOR2_X1 U516 ( .A1(n448), .A2(n452), .ZN(n454) );
  XNOR2_X1 U517 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n583), .A2(n551), .ZN(n455) );
  XNOR2_X1 U520 ( .A(KEYINPUT45), .B(n455), .ZN(n456) );
  NAND2_X1 U521 ( .A1(n456), .A2(n574), .ZN(n457) );
  NOR2_X1 U522 ( .A1(n555), .A2(n457), .ZN(n458) );
  AND2_X1 U523 ( .A1(n500), .A2(n543), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(KEYINPUT54), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n462), .A2(n512), .ZN(n567) );
  NOR2_X1 U526 ( .A1(n463), .A2(n567), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n467), .A2(n502), .ZN(n468) );
  INV_X1 U528 ( .A(n563), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n469), .A2(n535), .ZN(n472) );
  INV_X1 U530 ( .A(G183GAT), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n448), .A2(n551), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT97), .B(n476), .Z(n495) );
  NAND2_X1 U535 ( .A1(n477), .A2(n495), .ZN(n485) );
  NOR2_X1 U536 ( .A1(n512), .A2(n485), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT98), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NOR2_X1 U540 ( .A1(n514), .A2(n485), .ZN(n481) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n526), .A2(n485), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n484), .Z(G1326GAT) );
  NOR2_X1 U546 ( .A1(n520), .A2(n485), .ZN(n486) );
  XOR2_X1 U547 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  NOR2_X1 U548 ( .A1(n512), .A2(n490), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n514), .A2(n490), .ZN(n489) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  NOR2_X1 U553 ( .A1(n526), .A2(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  INV_X1 U558 ( .A(n512), .ZN(n497) );
  NAND2_X1 U559 ( .A1(n558), .A2(n541), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(KEYINPUT103), .ZN(n510) );
  NAND2_X1 U561 ( .A1(n510), .A2(n495), .ZN(n496) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n496), .Z(n506) );
  NAND2_X1 U563 ( .A1(n497), .A2(n506), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n500), .A2(n506), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n501), .ZN(G1333GAT) );
  XOR2_X1 U567 ( .A(G71GAT), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U568 ( .A1(n502), .A2(n506), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n508) );
  NAND2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n519) );
  NOR2_X1 U575 ( .A1(n512), .A2(n519), .ZN(n513) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n519), .ZN(n516) );
  XNOR2_X1 U578 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n519), .ZN(n518) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n543), .A2(n524), .ZN(n525) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n538), .A2(n555), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U592 ( .A1(n538), .A2(n558), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT112), .Z(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n533) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n537) );
  INV_X1 U599 ( .A(n538), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(n537), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U603 ( .A1(n538), .A2(n448), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT117), .Z(n547) );
  NOR2_X1 U606 ( .A1(n568), .A2(n542), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(n545), .Z(n553) );
  NAND2_X1 U609 ( .A1(n449), .A2(n553), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U612 ( .A1(n553), .A2(n558), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  INV_X1 U615 ( .A(n551), .ZN(n578) );
  NAND2_X1 U616 ( .A1(n553), .A2(n578), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n448), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U624 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .Z(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n448), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n570) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n577), .A2(n449), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(n571), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n577), .ZN(n582) );
  OR2_X1 U641 ( .A1(n582), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

