//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT88), .B(G29gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G36gat), .ZN(new_n204));
  OR3_X1    g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT87), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n204), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT15), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT89), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n212), .A2(new_n216), .A3(KEYINPUT15), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n207), .B1(new_n208), .B2(KEYINPUT90), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n219), .B(new_n204), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n213), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n219), .A2(new_n204), .ZN(new_n227));
  OAI221_X1 g026(.A(new_n227), .B1(new_n221), .B2(new_n222), .C1(new_n215), .C2(new_n217), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT17), .A3(new_n213), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n230), .A2(G1gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n230), .B(KEYINPUT91), .C1(new_n231), .C2(G1gat), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT92), .B(G8gat), .Z(new_n237));
  NAND4_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G8gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n241), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n202), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(G169gat), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT94), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n242), .A2(new_n228), .A3(new_n256), .A4(new_n213), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT94), .B1(new_n224), .B2(new_n241), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n245), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n244), .B(KEYINPUT13), .Z(new_n260));
  AOI22_X1  g059(.A1(new_n246), .A2(new_n247), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n244), .A4(new_n245), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n261), .B(new_n262), .C1(new_n248), .C2(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT96), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n264), .A2(KEYINPUT96), .A3(new_n265), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G141gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G148gat), .ZN(new_n272));
  INV_X1    g071(.A(G148gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G141gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT2), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n275), .A2(new_n276), .B1(G155gat), .B2(G162gat), .ZN(new_n277));
  INV_X1    g076(.A(G155gat), .ZN(new_n278));
  INV_X1    g077(.A(G162gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT72), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n272), .A2(new_n274), .B1(KEYINPUT2), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n283), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n284), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT73), .B1(new_n284), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n284), .A2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n282), .ZN(new_n296));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(G113gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(G120gat), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(G120gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT66), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n298), .ZN(new_n309));
  INV_X1    g108(.A(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n296), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n302), .A2(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n314), .A3(new_n282), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n292), .A2(new_n293), .B1(new_n281), .B2(new_n277), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT4), .A3(new_n314), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n313), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n313), .A2(new_n323), .A3(new_n317), .A4(new_n319), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT75), .B1(new_n325), .B2(KEYINPUT5), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n288), .A2(new_n312), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n329));
  INV_X1    g128(.A(new_n323), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n288), .A2(new_n331), .A3(new_n312), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n325), .A2(KEYINPUT5), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n334), .B1(new_n326), .B2(new_n324), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT6), .B1(new_n343), .B2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n341), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT76), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G226gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT23), .ZN(new_n369));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n359), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n375));
  AND3_X1   g174(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT24), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT65), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(G183gat), .B2(G190gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n381), .A3(new_n363), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n375), .B(KEYINPUT25), .C1(new_n378), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT27), .B(G183gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n365), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(KEYINPUT28), .A3(new_n365), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n368), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n360), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n374), .A2(new_n383), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n358), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n383), .A2(new_n374), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n389), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n357), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G197gat), .B(G204gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT22), .ZN(new_n403));
  INV_X1    g202(.A(G211gat), .ZN(new_n404));
  INV_X1    g203(.A(G218gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n402), .A3(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n400), .A3(new_n415), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n357), .B1(new_n399), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n395), .A2(new_n358), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n421), .B2(new_n412), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n354), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n412), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT71), .B1(new_n401), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(new_n414), .A3(new_n416), .A4(new_n353), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n417), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n425), .A4(new_n353), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n350), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n296), .A2(new_n418), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(new_n413), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n288), .A2(new_n418), .A3(new_n412), .ZN(new_n436));
  NAND2_X1  g235(.A1(G228gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n289), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n418), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT77), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n412), .A2(KEYINPUT77), .A3(new_n418), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n295), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n444), .A2(new_n288), .B1(new_n434), .B2(new_n424), .ZN(new_n445));
  OAI221_X1 g244(.A(new_n433), .B1(new_n435), .B2(new_n439), .C1(new_n445), .C2(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT31), .B(G50gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n288), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n424), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n438), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n439), .B1(new_n413), .B2(new_n434), .ZN(new_n455));
  OAI21_X1  g254(.A(G22gat), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n448), .A2(new_n451), .B1(new_n446), .B2(new_n456), .ZN(new_n457));
  AND4_X1   g256(.A1(KEYINPUT78), .A2(new_n446), .A3(new_n456), .A4(new_n451), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n399), .B2(new_n312), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n395), .A2(KEYINPUT67), .A3(new_n314), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n399), .A2(new_n312), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G15gat), .B(G43gat), .Z(new_n472));
  XNOR2_X1  g271(.A(G71gat), .B(G99gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n474), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n468), .B(KEYINPUT32), .C1(new_n470), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n465), .A2(new_n467), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n479), .B(KEYINPUT34), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n475), .A3(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT68), .B1(new_n478), .B2(new_n481), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(new_n481), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT69), .B1(new_n491), .B2(KEYINPUT36), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n460), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n341), .B1(new_n343), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n327), .A2(new_n498), .A3(new_n335), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n344), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n342), .ZN(new_n502));
  INV_X1    g301(.A(new_n426), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n423), .B1(new_n504), .B2(new_n353), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n401), .B2(new_n412), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n421), .A2(new_n413), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT38), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n502), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT82), .A4(new_n509), .ZN(new_n513));
  INV_X1    g312(.A(new_n505), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n504), .B1(new_n428), .B2(new_n425), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT38), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n313), .A2(new_n317), .A3(new_n319), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n330), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n521), .A3(new_n330), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n329), .A2(new_n332), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n526), .B2(new_n323), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n340), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(KEYINPUT40), .A3(new_n340), .A4(new_n528), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n531), .B(new_n532), .C1(new_n500), .C2(new_n499), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n431), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n459), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n517), .A2(new_n540), .A3(KEYINPUT83), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT83), .B1(new_n517), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n497), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n485), .A2(new_n459), .A3(new_n486), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n350), .A2(new_n545), .A3(new_n431), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n544), .A3(KEYINPUT35), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n491), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n501), .A2(new_n502), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR4_X1   g352(.A1(new_n550), .A2(new_n551), .A3(new_n459), .A4(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n270), .B1(new_n543), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  NAND2_X1  g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(G57gat), .A2(G64gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(G57gat), .A2(G64gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT97), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(KEYINPUT98), .A3(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n559), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n564), .A2(new_n565), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n572), .A2(new_n576), .A3(new_n558), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G127gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n241), .B1(KEYINPUT21), .B2(new_n579), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT100), .Z(new_n586));
  AND2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n584), .A2(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n278), .ZN(new_n591));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  NOR2_X1   g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n587), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT103), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(G92gat), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G99gat), .ZN(new_n609));
  INV_X1    g408(.A(G106gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT8), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n603), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G99gat), .B(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n603), .A2(new_n608), .A3(new_n613), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT101), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n224), .A2(new_n618), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n229), .A2(new_n617), .ZN(new_n623));
  INV_X1    g422(.A(new_n226), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT102), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n626), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n622), .B(new_n632), .C1(new_n623), .C2(new_n624), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n627), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n627), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n597), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n578), .A2(new_n617), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n575), .A2(new_n577), .A3(new_n615), .A4(new_n616), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g442(.A1(new_n575), .A2(new_n577), .A3(new_n615), .A4(new_n616), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n640), .B2(new_n642), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT104), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n647), .B(KEYINPUT105), .Z(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n643), .B2(new_n645), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n653), .B1(new_n658), .B2(new_n649), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n638), .A2(new_n639), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n594), .A2(new_n596), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n636), .ZN(new_n663));
  INV_X1    g462(.A(new_n660), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT106), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n557), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n557), .A2(KEYINPUT107), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n350), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  AND3_X1   g474(.A1(new_n671), .A2(new_n539), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G8gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n671), .B2(new_n539), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  INV_X1    g479(.A(new_n671), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n681), .A2(G15gat), .A3(new_n490), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n681), .B2(new_n496), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n671), .A2(new_n459), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  NAND3_X1  g486(.A1(new_n597), .A2(new_n637), .A3(new_n660), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT108), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n557), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n350), .A2(new_n203), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n460), .A2(new_n496), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n517), .A2(new_n540), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT83), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n517), .A2(new_n540), .A3(KEYINPUT83), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n546), .A2(new_n544), .A3(KEYINPUT35), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n547), .A3(new_n554), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n694), .B(new_n637), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n543), .A2(new_n556), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n706), .A2(new_n694), .A3(KEYINPUT44), .A4(new_n637), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n662), .A2(new_n267), .A3(new_n664), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n203), .B1(new_n709), .B2(new_n350), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n693), .A2(KEYINPUT110), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1328gat));
  INV_X1    g514(.A(new_n690), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(G36gat), .A3(new_n538), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n709), .B2(new_n538), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1329gat));
  OAI21_X1  g519(.A(G43gat), .B1(new_n709), .B2(new_n496), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n490), .A2(G43gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n690), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n724), .A2(KEYINPUT111), .A3(KEYINPUT47), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT47), .B1(new_n724), .B2(KEYINPUT111), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(new_n459), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n716), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n459), .A2(G50gat), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n729), .A2(G50gat), .B1(new_n709), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g531(.A1(new_n706), .A2(new_n267), .A3(new_n638), .A4(new_n664), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n672), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g534(.A(new_n538), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT112), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT113), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  INV_X1    g540(.A(new_n496), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n490), .A2(G71gat), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n743), .A2(G71gat), .B1(new_n733), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n733), .A2(new_n459), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g548(.A1(new_n662), .A2(new_n266), .A3(new_n660), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n705), .A2(new_n707), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n350), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n662), .A2(new_n266), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n637), .B(new_n753), .C1(new_n700), .C2(new_n702), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n637), .A4(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n672), .A2(new_n602), .A3(new_n664), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NOR3_X1   g560(.A1(new_n538), .A2(G92gat), .A3(new_n660), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n705), .A2(new_n539), .A3(new_n707), .A4(new_n750), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n599), .A2(new_n601), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n756), .A2(KEYINPUT115), .A3(new_n757), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n770), .A3(new_n755), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n771), .A3(new_n762), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n766), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  AOI211_X1 g574(.A(KEYINPUT116), .B(new_n775), .C1(new_n772), .C2(new_n766), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n774), .B2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n751), .B2(new_n496), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n491), .A2(new_n609), .A3(new_n664), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n759), .B2(new_n779), .ZN(G1338gat));
  OAI21_X1  g579(.A(G106gat), .B1(new_n751), .B2(new_n728), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n728), .A2(G106gat), .A3(new_n660), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n769), .A2(new_n771), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n758), .B2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n261), .A2(new_n254), .A3(new_n262), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n259), .A2(new_n260), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n253), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n636), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT54), .B(new_n657), .C1(new_n643), .C2(new_n645), .ZN(new_n795));
  INV_X1    g594(.A(new_n653), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT117), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  INV_X1    g597(.A(new_n657), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n575), .A2(new_n577), .B1(new_n615), .B2(new_n616), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n644), .A2(new_n800), .A3(KEYINPUT10), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n642), .A2(new_n641), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n798), .B(new_n799), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n653), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n798), .B1(new_n646), .B2(new_n647), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n643), .A2(new_n645), .A3(new_n657), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n807), .B2(new_n808), .ZN(new_n813));
  AOI211_X1 g612(.A(KEYINPUT117), .B(new_n796), .C1(new_n658), .C2(new_n798), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n804), .B1(new_n803), .B2(new_n653), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT118), .B1(new_n816), .B2(new_n656), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  AOI211_X1 g617(.A(new_n818), .B(new_n655), .C1(new_n806), .C2(new_n813), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n794), .B(new_n811), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n793), .A2(new_n660), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n656), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n818), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(KEYINPUT118), .A3(new_n656), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n810), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n825), .B2(new_n266), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT119), .B(new_n820), .C1(new_n826), .C2(new_n637), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n266), .B(new_n811), .C1(new_n819), .C2(new_n817), .ZN(new_n829));
  INV_X1    g628(.A(new_n821), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n637), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n820), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n827), .A2(new_n597), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n638), .A2(new_n267), .A3(new_n660), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n459), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n672), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n487), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n539), .ZN(new_n839));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n266), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n837), .A2(new_n538), .A3(new_n491), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n270), .A2(new_n300), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  AOI21_X1  g642(.A(G120gat), .B1(new_n839), .B2(new_n664), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n660), .A2(new_n303), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n841), .B2(new_n845), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n841), .A2(G127gat), .A3(new_n662), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT120), .Z(new_n848));
  AOI21_X1  g647(.A(G127gat), .B1(new_n839), .B2(new_n662), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n538), .A2(new_n637), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT121), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n838), .A2(G134gat), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n841), .A2(new_n637), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G134gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n496), .A2(new_n672), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n539), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n835), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n459), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n822), .A2(new_n810), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n268), .B2(new_n269), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n637), .B1(new_n865), .B2(new_n830), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n597), .B1(new_n866), .B2(new_n832), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n863), .B1(new_n867), .B2(new_n835), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n270), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n728), .B1(new_n834), .B2(new_n835), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n860), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n271), .C1(new_n269), .C2(new_n268), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT125), .Z(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT122), .B(new_n860), .C1(new_n862), .C2(new_n868), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n266), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n880), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT123), .B1(new_n880), .B2(G141gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n873), .B(KEYINPUT124), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n876), .B1(new_n884), .B2(new_n874), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n661), .A2(new_n270), .A3(new_n665), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n867), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n459), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n863), .B1(new_n834), .B2(new_n835), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n860), .A2(new_n664), .ZN(new_n891));
  OAI21_X1  g690(.A(G148gat), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n879), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n660), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n273), .A2(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n872), .A2(new_n273), .A3(new_n664), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1345gat));
  OAI21_X1  g698(.A(G155gat), .B1(new_n894), .B2(new_n597), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n872), .A2(new_n278), .A3(new_n662), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n894), .B2(new_n636), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n859), .A2(new_n852), .A3(G162gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n871), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n672), .A2(new_n538), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n834), .B2(new_n835), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n545), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n266), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n908), .A2(new_n490), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n836), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(G169gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n270), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n914), .B2(new_n916), .ZN(G1348gat));
  INV_X1    g716(.A(new_n914), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n918), .B2(new_n660), .ZN(new_n919));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n920), .A3(new_n664), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n364), .B1(new_n914), .B2(new_n662), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n662), .A2(new_n384), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n911), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n918), .B2(new_n636), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n928), .B2(new_n927), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n910), .A2(G190gat), .A3(new_n636), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n742), .A2(new_n728), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n909), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n266), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n890), .A2(new_n742), .A3(new_n908), .ZN(new_n940));
  INV_X1    g739(.A(G197gat), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n270), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(G1352gat));
  INV_X1    g742(.A(new_n940), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n944), .B2(new_n660), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n937), .A2(G204gat), .A3(new_n660), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n938), .A2(new_n404), .A3(new_n662), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n908), .A2(new_n742), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n662), .B(new_n950), .C1(new_n888), .C2(new_n889), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(G211gat), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n405), .A3(new_n637), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n940), .A2(new_n637), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n962), .B2(new_n405), .ZN(G1355gat));
endmodule


