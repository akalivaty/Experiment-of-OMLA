//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1349, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1424, new_n1425;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NOR2_X1   g0008(.A1(G58), .A2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n205), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n208), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT64), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n218), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n242), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(new_n250), .A3(G13), .A4(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n202), .B1(new_n250), .B2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n258), .A4(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n214), .A2(KEYINPUT67), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT15), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G87), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT8), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n214), .A2(new_n266), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n279), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT69), .B1(new_n269), .B2(new_n273), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n257), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n252), .A2(new_n254), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n264), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G238), .A4(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(G232), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n292), .B(new_n294), .C1(new_n225), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n213), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n299), .A2(new_n300), .B1(new_n303), .B2(new_n250), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT65), .B(G45), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n301), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n250), .A2(G274), .ZN(new_n307));
  AOI22_X1  g0107(.A1(G244), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n288), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT73), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n298), .A2(new_n308), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n288), .A2(KEYINPUT73), .A3(new_n311), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n288), .A2(KEYINPUT71), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT72), .B(G200), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n298), .B2(new_n308), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G190), .B2(new_n315), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n264), .A2(new_n285), .A3(new_n324), .A4(new_n287), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n327), .B(KEYINPUT74), .Z(new_n328));
  NAND2_X1  g0128(.A1(new_n286), .A2(new_n218), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n269), .A2(G77), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n258), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n255), .A2(new_n258), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n250), .A2(G20), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G68), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n330), .A2(new_n334), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n299), .A2(new_n300), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n290), .A2(new_n291), .A3(G232), .A4(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT77), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n295), .A2(new_n344), .A3(G232), .A4(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n290), .A2(new_n291), .A3(G226), .A4(new_n293), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n341), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(G238), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT13), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n345), .B2(new_n343), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n352), .C1(new_n356), .C2(new_n341), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n357), .A3(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n358), .B2(G169), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n340), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n340), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n358), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n354), .B2(new_n357), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(G226), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n290), .A2(new_n291), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G77), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n290), .A2(new_n291), .A3(G223), .A4(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT66), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n295), .A2(new_n376), .A3(G222), .A4(new_n293), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n290), .A2(new_n291), .A3(G222), .A4(new_n293), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT66), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n371), .B1(new_n380), .B2(new_n341), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(G179), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n267), .A2(new_n268), .B1(new_n276), .B2(new_n278), .ZN(new_n383));
  INV_X1    g0183(.A(G150), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n201), .A2(new_n214), .B1(new_n280), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n257), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n255), .A2(G50), .A3(new_n258), .A4(new_n337), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n252), .A2(new_n243), .A3(new_n254), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n381), .A2(new_n310), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(new_n321), .ZN(new_n394));
  INV_X1    g0194(.A(new_n375), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n379), .A2(new_n377), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n341), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n371), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(G190), .B(new_n371), .C1(new_n380), .C2(new_n341), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n389), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT9), .A4(new_n388), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n393), .B1(new_n404), .B2(KEYINPUT75), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT10), .B1(new_n404), .B2(new_n393), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n393), .B(KEYINPUT10), .C1(new_n404), .C2(KEYINPUT75), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n392), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n328), .A2(new_n364), .A3(new_n370), .A4(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n279), .A2(new_n337), .ZN(new_n411));
  INV_X1    g0211(.A(new_n279), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n336), .A2(new_n411), .B1(new_n286), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n275), .A2(new_n218), .ZN(new_n415));
  OAI21_X1  g0215(.A(G20), .B1(new_n415), .B2(new_n209), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n281), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n289), .B2(G33), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n266), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(G20), .B1(new_n422), .B2(new_n290), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n218), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n420), .B2(new_n421), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT7), .B1(new_n427), .B2(G20), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n418), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n258), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT16), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT79), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n289), .A3(G33), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n434), .A3(new_n291), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n424), .B1(new_n435), .B2(new_n214), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n295), .A2(KEYINPUT7), .A3(G20), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n436), .A2(new_n218), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n431), .B1(new_n438), .B2(new_n418), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n414), .B1(new_n430), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  INV_X1    g0241(.A(G226), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n293), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n422), .A2(new_n290), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n293), .A2(G223), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n427), .A2(new_n446), .B1(G33), .B2(G87), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n427), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n297), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n306), .A2(new_n307), .ZN(new_n452));
  INV_X1    g0252(.A(G232), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n303), .A2(new_n250), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n341), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n366), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n450), .B2(new_n297), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(G200), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n440), .A2(new_n441), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(G200), .B1(new_n451), .B2(new_n457), .ZN(new_n463));
  AOI211_X1 g0263(.A(G190), .B(new_n456), .C1(new_n450), .C2(new_n297), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n266), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT78), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n290), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n424), .A3(new_n214), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n428), .A3(G68), .ZN(new_n470));
  INV_X1    g0270(.A(new_n418), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(KEYINPUT16), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n435), .A2(new_n214), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT7), .ZN(new_n475));
  INV_X1    g0275(.A(new_n437), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(G68), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT16), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n413), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT81), .B1(new_n465), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n462), .A2(new_n480), .A3(KEYINPUT17), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n439), .A2(new_n257), .A3(new_n472), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n413), .C1(new_n463), .C2(new_n464), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT82), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n451), .A2(G179), .A3(new_n457), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n310), .B2(new_n459), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT18), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n410), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n226), .A2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G257), .B2(G1698), .ZN(new_n496));
  INV_X1    g0296(.A(G303), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n468), .A2(new_n496), .B1(new_n497), .B2(new_n295), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n297), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n302), .A2(G1), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  AND2_X1   g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(G274), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT84), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT5), .B(G41), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(G274), .A4(new_n500), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n500), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(G270), .A3(new_n341), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(KEYINPUT88), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT88), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g0312(.A(G190), .B(new_n499), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n214), .C1(G33), .C2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n257), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g0319(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n252), .A2(new_n517), .A3(new_n254), .ZN(new_n522));
  OR2_X1    g0322(.A1(KEYINPUT89), .A2(KEYINPUT20), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n519), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n250), .A2(G33), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n335), .A2(new_n517), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n498), .A2(new_n297), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n508), .A2(new_n510), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT88), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n508), .A2(KEYINPUT88), .A3(new_n510), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n513), .B(new_n528), .C1(new_n534), .C2(new_n368), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT21), .ZN(new_n536));
  OAI21_X1  g0336(.A(G169), .B1(new_n524), .B2(new_n527), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n524), .A2(new_n527), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(G179), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n499), .B1(new_n511), .B2(new_n512), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(KEYINPUT21), .A3(new_n539), .A4(G169), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n535), .A2(new_n538), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n335), .A2(new_n526), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n225), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT25), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n255), .B2(G107), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n545), .A2(G107), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n220), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n422), .A2(new_n214), .A3(new_n290), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n220), .A2(G20), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n550), .B1(new_n372), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n214), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n225), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n266), .A2(G20), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n552), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT24), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT22), .B1(new_n295), .B2(new_n553), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n558), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n552), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT90), .B1(new_n570), .B2(new_n257), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT90), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n572), .B(new_n258), .C1(new_n562), .C2(new_n569), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n549), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n509), .A2(G264), .A3(new_n341), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(G257), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1698), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n427), .A2(new_n578), .B1(G33), .B2(G294), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n579), .B2(new_n341), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n504), .A2(new_n507), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n316), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n310), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n580), .B2(new_n581), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n427), .A2(new_n578), .ZN(new_n589));
  INV_X1    g0389(.A(G294), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n266), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n297), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(G190), .A3(new_n508), .A4(new_n575), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n549), .C1(new_n571), .C2(new_n573), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n500), .A2(new_n221), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n341), .B1(G45), .B2(new_n307), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G238), .A2(G1698), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n224), .B2(G1698), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n427), .A2(new_n599), .B1(G33), .B2(G116), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n600), .B2(new_n341), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n394), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n366), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n269), .A2(G97), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n214), .B1(new_n348), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n220), .A2(new_n515), .A3(new_n225), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n427), .A2(new_n214), .A3(G68), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n257), .ZN(new_n611));
  INV_X1    g0411(.A(new_n273), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n286), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n545), .A2(G87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n545), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n611), .B(new_n613), .C1(new_n612), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n601), .A2(G169), .ZN(new_n619));
  OAI211_X1 g0419(.A(G179), .B(new_n597), .C1(new_n600), .C2(new_n341), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n544), .A2(new_n587), .A3(new_n595), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n475), .A2(G107), .A3(new_n476), .ZN(new_n626));
  XNOR2_X1  g0426(.A(G97), .B(G107), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT6), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n628), .A2(new_n515), .A3(G107), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n258), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n255), .A2(G97), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n255), .A2(G97), .A3(new_n258), .A4(new_n525), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n625), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n638), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n628), .B2(new_n627), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n641), .A2(new_n214), .B1(new_n202), .B2(new_n280), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n436), .A2(new_n437), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(G107), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT86), .B(new_n640), .C1(new_n644), .C2(new_n258), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n224), .A2(G1698), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n290), .B(new_n646), .C1(new_n466), .C2(new_n467), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT4), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT83), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n422), .A2(new_n650), .A3(new_n290), .A4(new_n646), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n646), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n290), .A2(new_n291), .A3(G250), .A4(G1698), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n514), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n341), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n509), .A2(new_n341), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n657), .A2(KEYINPUT85), .A3(new_n577), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT85), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n297), .B1(new_n505), .B2(new_n500), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(G257), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n508), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(G169), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n649), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n650), .B1(new_n427), .B2(new_n646), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n655), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n297), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT85), .B1(new_n657), .B2(new_n577), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n660), .A2(new_n659), .A3(G257), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n581), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(G179), .A3(new_n670), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n639), .A2(new_n645), .B1(new_n663), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(G200), .B1(new_n656), .B2(new_n662), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n634), .A2(new_n638), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(G190), .A3(new_n670), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT87), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n639), .A2(new_n645), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n663), .A2(new_n671), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n494), .A2(new_n624), .A3(new_n684), .ZN(G372));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n367), .A2(new_n369), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(new_n319), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(new_n364), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n485), .B1(new_n483), .B2(KEYINPUT81), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n690), .A2(new_n462), .B1(new_n484), .B2(new_n485), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n686), .B(new_n492), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n688), .B2(new_n364), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n490), .B(KEYINPUT18), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT94), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT95), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n402), .A2(new_n403), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT75), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n400), .A4(new_n399), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n697), .A2(KEYINPUT76), .A3(new_n400), .A4(new_n399), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n393), .A2(new_n699), .B1(new_n700), .B2(KEYINPUT10), .ZN(new_n701));
  INV_X1    g0501(.A(new_n408), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n407), .A2(KEYINPUT95), .A3(new_n408), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n692), .A2(new_n695), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n391), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n616), .A2(new_n622), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n709), .B2(new_n680), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n619), .A2(new_n711), .A3(new_n620), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n619), .B2(new_n620), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n618), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n674), .B1(new_n663), .B2(new_n671), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT26), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n714), .A3(new_n616), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n672), .A2(new_n676), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n714), .A2(new_n616), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n595), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n538), .A2(new_n542), .A3(new_n540), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n549), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n568), .B1(new_n567), .B2(new_n552), .ZN(new_n725));
  AND4_X1   g0525(.A1(new_n568), .A2(new_n552), .A3(new_n555), .A4(new_n560), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n257), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n572), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n257), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n730), .A2(KEYINPUT92), .A3(new_n585), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT92), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n574), .B2(new_n586), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n723), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT93), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT92), .B1(new_n730), .B2(new_n585), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n574), .A2(new_n732), .A3(new_n586), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n722), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n718), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n708), .B1(new_n494), .B2(new_n741), .ZN(G369));
  OAI21_X1  g0542(.A(new_n595), .B1(new_n730), .B2(new_n585), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n250), .A2(new_n214), .A3(G13), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT27), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT27), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(G213), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G343), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n730), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT96), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n574), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT96), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n587), .A2(new_n753), .A3(new_n754), .A4(new_n595), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n587), .A2(new_n750), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n528), .A2(new_n750), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n722), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n543), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n737), .A2(new_n738), .A3(new_n750), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n723), .A2(new_n749), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n752), .A2(new_n755), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(G399));
  INV_X1    g0569(.A(new_n206), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G41), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n607), .A2(G116), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n772), .A2(G1), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n211), .B2(new_n772), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT97), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n741), .B2(new_n749), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n716), .B1(new_n720), .B2(new_n715), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n709), .A2(new_n680), .A3(KEYINPUT26), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n714), .B(KEYINPUT98), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n595), .A2(new_n616), .A3(new_n714), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n680), .A2(new_n682), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n587), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n722), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n749), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT29), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n778), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n734), .A2(new_n735), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n740), .A3(new_n785), .ZN(new_n793));
  INV_X1    g0593(.A(new_n718), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n749), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n789), .B1(new_n795), .B2(new_n777), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G330), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT30), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n580), .A2(new_n601), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(new_n667), .A3(new_n670), .ZN(new_n801));
  OAI211_X1 g0601(.A(G179), .B(new_n499), .C1(new_n511), .C2(new_n512), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n601), .A2(new_n316), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n582), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n805), .B(new_n541), .C1(new_n656), .C2(new_n662), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n801), .A2(new_n802), .A3(new_n799), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n749), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT31), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(KEYINPUT31), .B(new_n749), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n743), .A2(new_n543), .A3(new_n709), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n814), .A2(new_n677), .A3(new_n683), .A4(new_n750), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n798), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n776), .B1(new_n817), .B2(G1), .ZN(G364));
  AND2_X1   g0618(.A1(new_n214), .A2(G13), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n250), .B1(new_n819), .B2(G45), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n772), .A2(KEYINPUT99), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT99), .ZN(new_n822));
  INV_X1    g0622(.A(new_n820), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n771), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n764), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(G330), .B2(new_n762), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n213), .B1(G20), .B2(new_n310), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n427), .A2(new_n770), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n212), .A2(new_n305), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n248), .C2(new_n302), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n770), .A2(new_n372), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G355), .B1(new_n517), .B2(new_n770), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n366), .A2(G179), .A3(G200), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n214), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n515), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n214), .A2(G179), .ZN(new_n844));
  NOR2_X1   g0644(.A1(G190), .A2(G200), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n843), .B1(KEYINPUT32), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n214), .A2(new_n316), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n845), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n295), .B1(new_n852), .B2(new_n202), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(G190), .A3(new_n368), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(G58), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n394), .A2(new_n844), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(G190), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n225), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n366), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n857), .B(new_n861), .C1(G87), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n851), .A2(G200), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n366), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(G190), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G50), .A2(new_n865), .B1(new_n866), .B2(G68), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n863), .B(new_n867), .C1(KEYINPUT32), .C2(new_n849), .ZN(new_n868));
  INV_X1    g0668(.A(G322), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n854), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G311), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n372), .B1(new_n852), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n846), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n870), .B(new_n872), .C1(G329), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n862), .A2(G303), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G283), .B2(new_n859), .ZN(new_n877));
  INV_X1    g0677(.A(new_n842), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G294), .A2(new_n878), .B1(new_n865), .B2(G326), .ZN(new_n879));
  INV_X1    g0679(.A(new_n866), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT33), .B(G317), .Z(new_n881));
  OAI211_X1 g0681(.A(new_n877), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n868), .A2(new_n882), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n825), .B(new_n840), .C1(new_n883), .C2(new_n832), .ZN(new_n884));
  INV_X1    g0684(.A(new_n831), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n762), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n828), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G396));
  OAI21_X1  g0688(.A(new_n785), .B1(new_n739), .B2(KEYINPUT93), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n735), .B(new_n722), .C1(new_n737), .C2(new_n738), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n794), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n750), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n318), .A2(new_n317), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT73), .B1(new_n288), .B2(new_n311), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n326), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n288), .A2(new_n749), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n897), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n320), .A2(new_n325), .A3(new_n323), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n319), .B(new_n899), .C1(new_n893), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n891), .A2(new_n750), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n813), .A2(new_n815), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n826), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n816), .A3(new_n905), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n852), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n855), .A2(G143), .B1(new_n912), .B2(G159), .ZN(new_n913));
  INV_X1    g0713(.A(G137), .ZN(new_n914));
  INV_X1    g0714(.A(new_n865), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n913), .B1(new_n880), .B2(new_n384), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT34), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n859), .A2(G68), .ZN(new_n918));
  INV_X1    g0718(.A(new_n862), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n243), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G132), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n427), .B1(new_n923), .B2(new_n846), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(KEYINPUT101), .B1(G58), .B2(new_n878), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(KEYINPUT101), .B2(new_n924), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n843), .B1(G303), .B2(new_n865), .ZN(new_n927));
  INV_X1    g0727(.A(G283), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n880), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n854), .A2(new_n590), .B1(new_n852), .B2(new_n517), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n295), .B(new_n930), .C1(G311), .C2(new_n873), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n862), .A2(G107), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n859), .A2(G87), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n922), .A2(new_n926), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n832), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n832), .A2(new_n829), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n825), .B1(new_n202), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n829), .B2(new_n902), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n911), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(G384));
  OR2_X1    g0742(.A1(new_n632), .A2(KEYINPUT35), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n632), .A2(KEYINPUT35), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(G116), .A3(new_n215), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  OR3_X1    g0746(.A1(new_n211), .A2(new_n202), .A3(new_n415), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n244), .B(KEYINPUT103), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n250), .B(G13), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT38), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n429), .A2(KEYINPUT16), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n413), .B1(new_n952), .B2(new_n473), .ZN(new_n953));
  INV_X1    g0753(.A(new_n747), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n487), .B2(new_n492), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT37), .B1(new_n479), .B2(new_n489), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n440), .A2(new_n441), .A3(new_n460), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n480), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT104), .B1(new_n479), .B2(new_n954), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n961), .B(new_n747), .C1(new_n482), .C2(new_n413), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n953), .B1(new_n489), .B2(new_n954), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n480), .A2(new_n964), .A3(new_n958), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n959), .A2(new_n963), .B1(new_n965), .B2(KEYINPUT37), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n951), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n959), .A2(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(KEYINPUT37), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n955), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n691), .B2(new_n694), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT38), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n340), .A2(new_n749), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n370), .A2(new_n364), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n358), .A2(G169), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT14), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n361), .A3(new_n360), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n340), .B(new_n749), .C1(new_n687), .C2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n902), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n624), .A2(new_n684), .A3(new_n749), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n811), .A2(new_n812), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n974), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n963), .B1(new_n487), .B2(new_n492), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n490), .B(new_n483), .C1(new_n960), .C2(new_n962), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n963), .A2(new_n959), .B1(new_n991), .B2(KEYINPUT37), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n973), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n981), .B(KEYINPUT40), .C1(new_n982), .C2(new_n983), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n986), .A2(new_n988), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n494), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n997), .A2(new_n998), .A3(new_n907), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n907), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n798), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n319), .A2(new_n749), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n905), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n976), .A2(new_n980), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n974), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT39), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n956), .A2(new_n966), .A3(new_n951), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n989), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n991), .A2(KEYINPUT37), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n968), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n960), .A2(new_n962), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n691), .B2(new_n694), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1009), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1007), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n979), .A2(new_n340), .A3(new_n750), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n967), .A2(new_n973), .A3(KEYINPUT39), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n694), .A2(new_n747), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1006), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n707), .B1(new_n797), .B2(new_n998), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1001), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n250), .B2(new_n819), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1001), .A2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n950), .B1(new_n1025), .B2(new_n1026), .ZN(G367));
  NAND2_X1  g0827(.A1(new_n615), .A2(new_n749), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n720), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT107), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n714), .A2(new_n1028), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n720), .A2(KEYINPUT107), .A3(new_n1028), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT108), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1036), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT43), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1035), .A2(new_n1039), .A3(new_n1037), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n719), .B1(new_n674), .B2(new_n750), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n715), .A2(new_n749), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n680), .B1(new_n1046), .B2(new_n587), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n750), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n768), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT42), .B1(new_n1049), .B2(new_n1045), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT42), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1046), .A2(new_n768), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1040), .A2(new_n1042), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT109), .B1(new_n1053), .B2(new_n1042), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT109), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1056), .A2(new_n1057), .A3(new_n1041), .A4(new_n1048), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n765), .A2(new_n1046), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n771), .B(KEYINPUT41), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n768), .A2(new_n766), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n1046), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT44), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(KEYINPUT44), .A3(new_n1046), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT45), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1063), .B2(new_n1046), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n766), .A4(new_n1045), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1068), .A2(new_n765), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n765), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n892), .A2(KEYINPUT97), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n789), .A2(new_n1076), .B1(new_n778), .B2(new_n790), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT110), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n757), .B(new_n767), .C1(new_n752), .C2(new_n755), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n764), .B1(new_n1079), .B2(new_n1049), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n763), .B(new_n768), .C1(new_n759), .C2(new_n767), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1078), .A3(new_n908), .A4(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n791), .A2(new_n796), .A3(new_n1082), .A4(new_n908), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT110), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1075), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1062), .B1(new_n1086), .B2(new_n817), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1061), .B1(new_n1087), .B2(new_n823), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1038), .A2(new_n831), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n238), .A2(new_n770), .A3(new_n427), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n833), .B1(new_n206), .B2(new_n612), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n826), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n862), .A2(G116), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT46), .Z(new_n1094));
  INV_X1    g0894(.A(G317), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n854), .A2(new_n497), .B1(new_n846), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G283), .B2(new_n912), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n859), .A2(G97), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n427), .B1(new_n866), .B2(G294), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G107), .A2(new_n878), .B1(new_n865), .B2(G311), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n842), .A2(new_n218), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G143), .B2(new_n865), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n847), .B2(new_n880), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n854), .A2(new_n384), .B1(new_n852), .B2(new_n243), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n372), .B(new_n1105), .C1(G137), .C2(new_n873), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n859), .A2(G77), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n862), .A2(G58), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1094), .A2(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT47), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1092), .B1(new_n1111), .B2(new_n832), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1088), .A2(new_n1113), .ZN(G387));
  NAND2_X1  g0914(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n771), .C1(new_n817), .C2(new_n1082), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n756), .A2(new_n758), .A3(new_n831), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n835), .B1(new_n234), .B2(new_n305), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n838), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n773), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n412), .B2(G50), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n279), .A2(new_n1121), .A3(new_n243), .ZN(new_n1124));
  AOI21_X1  g0924(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n773), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1120), .A2(new_n1126), .B1(new_n225), .B2(new_n770), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n826), .B1(new_n1127), .B2(new_n834), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G68), .A2(new_n912), .B1(new_n873), .B2(G150), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n243), .B2(new_n854), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G97), .B2(new_n859), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n847), .A2(new_n915), .B1(new_n880), .B2(new_n412), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n842), .A2(new_n612), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1132), .A2(new_n468), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n862), .A2(G77), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n880), .A2(new_n871), .B1(new_n915), .B2(new_n869), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1137), .A2(KEYINPUT112), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(KEYINPUT112), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n855), .A2(G317), .B1(new_n912), .B2(G303), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT48), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n919), .A2(new_n590), .B1(new_n928), .B2(new_n842), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(KEYINPUT49), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n427), .B1(G326), .B2(new_n873), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n517), .C2(new_n860), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT49), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1136), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1128), .B1(new_n1150), .B2(new_n832), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1082), .A2(new_n823), .B1(new_n1117), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1116), .A2(new_n1152), .ZN(G393));
  AOI21_X1  g0953(.A(KEYINPUT44), .B1(new_n1063), .B2(new_n1046), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1067), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1072), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n764), .A3(new_n759), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT113), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1068), .A2(new_n765), .A3(new_n1072), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT113), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n823), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n873), .A2(G143), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n919), .B2(new_n218), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT114), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT114), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1165), .A2(new_n427), .A3(new_n933), .A4(new_n1166), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT115), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n842), .A2(new_n202), .B1(new_n412), .B2(new_n852), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G150), .A2(new_n865), .B1(new_n855), .B2(G159), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT51), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G50), .C2(new_n866), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT116), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n372), .B1(new_n846), .B2(new_n869), .C1(new_n590), .C2(new_n852), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1175), .B(new_n861), .C1(G283), .C2(new_n862), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n915), .A2(new_n1095), .B1(new_n871), .B2(new_n854), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT52), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n880), .A2(new_n497), .B1(new_n517), .B2(new_n842), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT117), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1174), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1168), .A2(KEYINPUT116), .A3(new_n1173), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n832), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n242), .A2(new_n835), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n834), .B1(G97), .B2(new_n770), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n825), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(new_n1045), .C2(new_n885), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1086), .A2(new_n771), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1075), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1162), .B(new_n1188), .C1(new_n1189), .C2(new_n1190), .ZN(G390));
  AND3_X1   g0991(.A1(new_n967), .A2(KEYINPUT39), .A3(new_n973), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT39), .B1(new_n993), .B2(new_n973), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n829), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n937), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n826), .B1(new_n279), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n915), .A2(new_n1197), .B1(new_n923), .B2(new_n854), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT118), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n880), .A2(new_n914), .B1(new_n847), .B2(new_n842), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n372), .B1(new_n873), .B2(G125), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT54), .B(G143), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n852), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1199), .B(new_n1204), .C1(new_n243), .C2(new_n860), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n862), .A2(G150), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT53), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G77), .A2(new_n878), .B1(new_n865), .B2(G283), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n225), .B2(new_n880), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n862), .A2(G87), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n295), .B1(new_n912), .B2(G97), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n855), .A2(G116), .B1(new_n873), .B2(G294), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n918), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1205), .A2(new_n1207), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1196), .B1(new_n1214), .B2(new_n832), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1005), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n905), .B2(new_n1003), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1218), .A2(new_n1017), .B1(new_n1193), .B2(new_n1192), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1002), .B1(new_n788), .B2(new_n904), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1016), .B(new_n994), .C1(new_n1220), .C2(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n816), .A2(new_n904), .A3(new_n1005), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n816), .A2(new_n904), .A3(new_n1005), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1219), .A2(new_n1225), .A3(new_n1221), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1216), .B1(new_n1227), .B2(new_n820), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n494), .A2(new_n908), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n707), .B(new_n1229), .C1(new_n797), .C2(new_n998), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1005), .B1(new_n816), .B2(new_n904), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1004), .B1(new_n1223), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1217), .B1(new_n908), .B2(new_n902), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1225), .A3(new_n1220), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1224), .A2(new_n1230), .A3(new_n1226), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1229), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1022), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n772), .B1(new_n1227), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1228), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G378));
  NAND2_X1  g1041(.A1(new_n389), .A2(new_n954), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT55), .Z(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT120), .B1(new_n705), .B2(new_n391), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT120), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1245), .B(new_n392), .C1(new_n703), .C2(new_n704), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n407), .A2(KEYINPUT95), .A3(new_n408), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT95), .B1(new_n407), .B2(new_n408), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n391), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1245), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1243), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n705), .A2(KEYINPUT120), .A3(new_n391), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1247), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1248), .B1(new_n1247), .B2(new_n1255), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n829), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n859), .A2(G58), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G41), .B1(new_n912), .B2(new_n273), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n855), .A2(G107), .B1(new_n873), .B2(G283), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1135), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n880), .A2(new_n515), .B1(new_n915), .B2(new_n517), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1263), .A2(new_n427), .A3(new_n1102), .A4(new_n1264), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT58), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(KEYINPUT58), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G41), .B1(new_n427), .B2(G33), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1267), .C1(G50), .C2(new_n1268), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n854), .A2(new_n1197), .B1(new_n852), .B2(new_n914), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G132), .B2(new_n866), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G150), .A2(new_n878), .B1(new_n865), .B2(G125), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1271), .B(new_n1272), .C1(new_n919), .C2(new_n1202), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT59), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n859), .A2(G159), .ZN(new_n1275));
  AOI211_X1 g1075(.A(G33), .B(G41), .C1(new_n873), .C2(G124), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1273), .A2(KEYINPUT59), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n832), .B1(new_n1269), .B2(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT119), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n937), .A2(new_n243), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1259), .A2(new_n826), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1248), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1244), .A2(new_n1246), .A3(new_n1243), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1253), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1247), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n997), .A3(G330), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n996), .A2(new_n994), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n984), .B1(new_n973), .B2(new_n967), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1291), .B(G330), .C1(new_n1292), .C2(new_n987), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1258), .A2(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1290), .A2(new_n1294), .A3(new_n1021), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1021), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1283), .B1(new_n1297), .B2(new_n820), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1237), .B(new_n708), .C1(new_n1077), .C2(new_n494), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1219), .A2(new_n1225), .A3(new_n1221), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1225), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1303), .B2(new_n1235), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT57), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n771), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1236), .A2(new_n1230), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1021), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1289), .B1(G330), .B2(new_n997), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1258), .A2(new_n1293), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1290), .A2(new_n1294), .A3(new_n1021), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT57), .B1(new_n1307), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1299), .B1(new_n1306), .B2(new_n1314), .ZN(G375));
  NAND2_X1  g1115(.A1(new_n1217), .A2(new_n829), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n826), .B1(G68), .B2(new_n1195), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n866), .A2(G116), .B1(new_n912), .B2(G107), .ZN(new_n1318));
  XOR2_X1   g1118(.A(new_n1318), .B(KEYINPUT122), .Z(new_n1319));
  AOI21_X1  g1119(.A(new_n1133), .B1(G294), .B2(new_n865), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n862), .A2(G97), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n372), .B1(new_n854), .B2(new_n928), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(G303), .B2(new_n873), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1107), .A2(new_n1320), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n468), .B1(new_n865), .B2(G132), .ZN(new_n1325));
  OAI221_X1 g1125(.A(new_n1325), .B1(new_n243), .B2(new_n842), .C1(new_n880), .C2(new_n1202), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n862), .A2(G159), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n912), .A2(G150), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n855), .A2(G137), .B1(new_n873), .B2(G128), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1260), .A2(new_n1327), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  OAI22_X1  g1130(.A1(new_n1319), .A2(new_n1324), .B1(new_n1326), .B2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1317), .B1(new_n1331), .B2(new_n832), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1235), .A2(new_n823), .B1(new_n1316), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1062), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1238), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1235), .B1(new_n1022), .B2(new_n1237), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(G381));
  NOR4_X1   g1137(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1338));
  INV_X1    g1138(.A(G390), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(new_n1088), .A3(new_n1113), .A4(new_n1339), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1340), .A2(KEYINPUT123), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT57), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1342), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n772), .B1(new_n1343), .B2(new_n1307), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1304), .B2(new_n1297), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1298), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1340), .A2(KEYINPUT123), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1341), .A2(new_n1240), .A3(new_n1346), .A4(new_n1347), .ZN(G407));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1240), .ZN(new_n1349));
  OAI211_X1 g1149(.A(G407), .B(G213), .C1(G343), .C2(new_n1349), .ZN(G409));
  AOI21_X1  g1150(.A(new_n1336), .B1(KEYINPUT60), .B2(new_n1238), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1300), .A2(new_n1352), .A3(KEYINPUT60), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n771), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1333), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n941), .ZN(new_n1356));
  OAI211_X1 g1156(.A(G384), .B(new_n1333), .C1(new_n1351), .C2(new_n1354), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(G2897), .ZN(new_n1359));
  INV_X1    g1159(.A(G213), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1360), .A2(G343), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1358), .B1(new_n1359), .B2(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1359), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1356), .A2(new_n1357), .A3(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(KEYINPUT124), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT124), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1311), .A2(new_n1368), .A3(new_n1312), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1367), .A2(new_n1369), .A3(new_n823), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1307), .A2(new_n1334), .A3(new_n1313), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1240), .A2(new_n1283), .A3(new_n1370), .A4(new_n1371), .ZN(new_n1372));
  OAI211_X1 g1172(.A(new_n1362), .B(new_n1372), .C1(new_n1346), .C2(new_n1240), .ZN(new_n1373));
  AOI21_X1  g1173(.A(KEYINPUT61), .B1(new_n1366), .B2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1240), .B1(new_n1375), .B2(new_n1299), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1227), .A2(new_n1238), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(new_n1236), .A3(new_n771), .ZN(new_n1379));
  AOI22_X1  g1179(.A1(new_n1303), .A2(new_n823), .B1(new_n1194), .B2(new_n1215), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1379), .A2(new_n1380), .A3(new_n1283), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1362), .B1(new_n1377), .B2(new_n1381), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1376), .A2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1358), .ZN(new_n1384));
  AND3_X1   g1184(.A1(new_n1383), .A2(KEYINPUT62), .A3(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT62), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1374), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1387));
  XNOR2_X1  g1187(.A(G393), .B(G396), .ZN(new_n1388));
  AND3_X1   g1188(.A1(new_n1088), .A2(new_n1113), .A3(G390), .ZN(new_n1389));
  AOI21_X1  g1189(.A(G390), .B1(new_n1088), .B2(new_n1113), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1388), .B1(new_n1389), .B2(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(G387), .A2(new_n1339), .ZN(new_n1392));
  XNOR2_X1  g1192(.A(G393), .B(new_n887), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1088), .A2(new_n1113), .A3(G390), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1392), .A2(new_n1393), .A3(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1391), .A2(new_n1395), .ZN(new_n1396));
  XNOR2_X1  g1196(.A(new_n1396), .B(KEYINPUT127), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1387), .A2(new_n1397), .ZN(new_n1398));
  AND2_X1   g1198(.A1(new_n1391), .A2(new_n1395), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT61), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(G375), .A2(G378), .ZN(new_n1401));
  AOI21_X1  g1201(.A(new_n820), .B1(new_n1313), .B2(KEYINPUT124), .ZN(new_n1402));
  AOI22_X1  g1202(.A1(new_n1236), .A2(new_n1230), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1403));
  AOI22_X1  g1203(.A1(new_n1402), .A2(new_n1369), .B1(new_n1403), .B2(new_n1334), .ZN(new_n1404));
  AND3_X1   g1204(.A1(new_n1379), .A2(new_n1380), .A3(new_n1283), .ZN(new_n1405));
  AOI21_X1  g1205(.A(new_n1361), .B1(new_n1404), .B2(new_n1405), .ZN(new_n1406));
  AND3_X1   g1206(.A1(new_n1356), .A2(KEYINPUT63), .A3(new_n1357), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1401), .A2(new_n1406), .A3(new_n1407), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1399), .A2(new_n1400), .A3(new_n1408), .ZN(new_n1409));
  AOI21_X1  g1209(.A(KEYINPUT63), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1410));
  NOR2_X1   g1210(.A1(new_n1409), .A2(new_n1410), .ZN(new_n1411));
  OAI21_X1  g1211(.A(KEYINPUT125), .B1(new_n1376), .B2(new_n1382), .ZN(new_n1412));
  INV_X1    g1212(.A(KEYINPUT125), .ZN(new_n1413));
  NAND3_X1  g1213(.A1(new_n1401), .A2(new_n1406), .A3(new_n1413), .ZN(new_n1414));
  NAND3_X1  g1214(.A1(new_n1412), .A2(new_n1414), .A3(new_n1366), .ZN(new_n1415));
  AOI21_X1  g1215(.A(KEYINPUT126), .B1(new_n1411), .B2(new_n1415), .ZN(new_n1416));
  INV_X1    g1216(.A(KEYINPUT63), .ZN(new_n1417));
  OAI21_X1  g1217(.A(new_n1417), .B1(new_n1373), .B2(new_n1358), .ZN(new_n1418));
  NAND4_X1  g1218(.A1(new_n1418), .A2(new_n1400), .A3(new_n1399), .A4(new_n1408), .ZN(new_n1419));
  AND3_X1   g1219(.A1(new_n1412), .A2(new_n1414), .A3(new_n1366), .ZN(new_n1420));
  INV_X1    g1220(.A(KEYINPUT126), .ZN(new_n1421));
  NOR3_X1   g1221(.A1(new_n1419), .A2(new_n1420), .A3(new_n1421), .ZN(new_n1422));
  OAI21_X1  g1222(.A(new_n1398), .B1(new_n1416), .B2(new_n1422), .ZN(G405));
  NAND2_X1  g1223(.A1(new_n1401), .A2(new_n1349), .ZN(new_n1424));
  XNOR2_X1  g1224(.A(new_n1424), .B(new_n1358), .ZN(new_n1425));
  XNOR2_X1  g1225(.A(new_n1425), .B(new_n1396), .ZN(G402));
endmodule


