

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n738), .A2(n737), .ZN(n741) );
  AND2_X1 U555 ( .A1(G137), .A2(n889), .ZN(n520) );
  XOR2_X1 U556 ( .A(KEYINPUT101), .B(n733), .Z(n521) );
  AND2_X1 U557 ( .A1(G1976), .A2(G288), .ZN(n522) );
  AND2_X1 U558 ( .A1(n965), .A2(n827), .ZN(n523) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n711) );
  INV_X1 U560 ( .A(KEYINPUT102), .ZN(n739) );
  XNOR2_X1 U561 ( .A(n739), .B(KEYINPUT31), .ZN(n740) );
  XNOR2_X1 U562 ( .A(n741), .B(n740), .ZN(n742) );
  BUF_X1 U563 ( .A(n710), .Z(n744) );
  NOR2_X1 U564 ( .A1(G1966), .A2(n774), .ZN(n756) );
  AND2_X1 U565 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U566 ( .A1(n699), .A2(n801), .ZN(n710) );
  INV_X1 U567 ( .A(G2104), .ZN(n525) );
  OR2_X1 U568 ( .A1(n814), .A2(n523), .ZN(n815) );
  NOR2_X2 U569 ( .A1(G2105), .A2(n525), .ZN(n888) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n652) );
  XNOR2_X1 U571 ( .A(n524), .B(KEYINPUT65), .ZN(n893) );
  AND2_X1 U572 ( .A1(n532), .A2(n531), .ZN(G160) );
  NAND2_X1 U573 ( .A1(n525), .A2(G2105), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G125), .A2(n893), .ZN(n532) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U576 ( .A1(n892), .A2(G113), .ZN(n528) );
  NAND2_X1 U577 ( .A1(G101), .A2(n888), .ZN(n526) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n529), .Z(n889) );
  NOR2_X1 U582 ( .A1(n530), .A2(n520), .ZN(n531) );
  XOR2_X1 U583 ( .A(G2446), .B(KEYINPUT106), .Z(n534) );
  XNOR2_X1 U584 ( .A(G2451), .B(G2430), .ZN(n533) );
  XNOR2_X1 U585 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U586 ( .A(n535), .B(G2427), .Z(n537) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U588 ( .A(n537), .B(n536), .ZN(n541) );
  XOR2_X1 U589 ( .A(G2443), .B(G2435), .Z(n539) );
  XNOR2_X1 U590 ( .A(G2438), .B(G2454), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U592 ( .A(n541), .B(n540), .Z(n542) );
  AND2_X1 U593 ( .A1(G14), .A2(n542), .ZN(G401) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U595 ( .A(G132), .ZN(G219) );
  INV_X1 U596 ( .A(G82), .ZN(G220) );
  INV_X1 U597 ( .A(G120), .ZN(G236) );
  INV_X1 U598 ( .A(G69), .ZN(G235) );
  INV_X1 U599 ( .A(G108), .ZN(G238) );
  INV_X1 U600 ( .A(G651), .ZN(n548) );
  NOR2_X1 U601 ( .A1(G543), .A2(n548), .ZN(n543) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n543), .Z(n651) );
  NAND2_X1 U603 ( .A1(G62), .A2(n651), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  NOR2_X1 U605 ( .A1(G651), .A2(n644), .ZN(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT64), .B(n544), .ZN(n653) );
  NAND2_X1 U607 ( .A1(G50), .A2(n653), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT84), .B(n547), .Z(n552) );
  NAND2_X1 U610 ( .A1(G88), .A2(n652), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n644), .A2(n548), .ZN(n658) );
  NAND2_X1 U612 ( .A1(G75), .A2(n658), .ZN(n549) );
  AND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(G303) );
  XOR2_X1 U615 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n554) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(G223) );
  INV_X1 U618 ( .A(G223), .ZN(n832) );
  NAND2_X1 U619 ( .A1(n832), .A2(G567), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U621 ( .A1(n651), .A2(G56), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT14), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G43), .A2(n653), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT70), .B(KEYINPUT12), .Z(n560) );
  NAND2_X1 U626 ( .A1(G81), .A2(n652), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n658), .A2(G68), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT71), .B(n561), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT73), .ZN(n974) );
  INV_X1 U635 ( .A(G860), .ZN(n628) );
  OR2_X1 U636 ( .A1(n974), .A2(n628), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G64), .A2(n651), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G52), .A2(n653), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G90), .A2(n652), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G77), .A2(n658), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT66), .B(n576), .Z(G301) );
  NAND2_X1 U646 ( .A1(G301), .A2(G868), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G79), .A2(n658), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n652), .A2(G92), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G54), .A2(n653), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n651), .A2(G66), .ZN(n579) );
  XOR2_X1 U652 ( .A(KEYINPUT74), .B(n579), .Z(n580) );
  NOR2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT15), .ZN(n861) );
  INV_X1 U656 ( .A(n861), .ZN(n977) );
  INV_X1 U657 ( .A(G868), .ZN(n669) );
  NAND2_X1 U658 ( .A1(n977), .A2(n669), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U660 ( .A1(n651), .A2(G65), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G78), .A2(n658), .ZN(n587) );
  XOR2_X1 U662 ( .A(KEYINPUT67), .B(n587), .Z(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n652), .A2(G91), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G53), .A2(n653), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n967) );
  XOR2_X1 U668 ( .A(n967), .B(KEYINPUT68), .Z(G299) );
  NAND2_X1 U669 ( .A1(n651), .A2(G63), .ZN(n594) );
  XOR2_X1 U670 ( .A(KEYINPUT77), .B(n594), .Z(n596) );
  NAND2_X1 U671 ( .A1(G51), .A2(n653), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n598) );
  XOR2_X1 U673 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n597) );
  XOR2_X1 U674 ( .A(n598), .B(n597), .Z(n606) );
  NAND2_X1 U675 ( .A1(n658), .A2(G76), .ZN(n599) );
  XOR2_X1 U676 ( .A(KEYINPUT76), .B(n599), .Z(n603) );
  NAND2_X1 U677 ( .A1(G89), .A2(n652), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT4), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT75), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U681 ( .A(KEYINPUT5), .B(n604), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n607), .B(KEYINPUT79), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U685 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U686 ( .A1(G299), .A2(G868), .ZN(n610) );
  NOR2_X1 U687 ( .A1(G286), .A2(n669), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n628), .A2(G559), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n611), .A2(n861), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U692 ( .A1(G559), .A2(n977), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n613), .A2(G868), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n974), .A2(n669), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U696 ( .A1(n892), .A2(G111), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n616), .B(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G99), .A2(n888), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT81), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G135), .A2(n889), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n893), .A2(G123), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT18), .B(n622), .Z(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n927) );
  XNOR2_X1 U706 ( .A(G2096), .B(n927), .ZN(n626) );
  INV_X1 U707 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U709 ( .A1(G559), .A2(n861), .ZN(n627) );
  XOR2_X1 U710 ( .A(n974), .B(n627), .Z(n666) );
  NAND2_X1 U711 ( .A1(n628), .A2(n666), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G93), .A2(n652), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G80), .A2(n658), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U715 ( .A(KEYINPUT82), .B(n631), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G67), .A2(n651), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G55), .A2(n653), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n668) );
  XOR2_X1 U720 ( .A(n636), .B(n668), .Z(G145) );
  INV_X1 U721 ( .A(G303), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G61), .A2(n651), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G48), .A2(n653), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n658), .A2(G73), .ZN(n639) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n652), .A2(G86), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U730 ( .A1(n644), .A2(G87), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G49), .A2(n653), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n651), .A2(n647), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n648) );
  XOR2_X1 U735 ( .A(KEYINPUT83), .B(n648), .Z(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G288) );
  AND2_X1 U737 ( .A1(n651), .A2(G60), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n652), .A2(G85), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G47), .A2(n653), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n658), .A2(G72), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(G290) );
  XNOR2_X1 U744 ( .A(KEYINPUT19), .B(n668), .ZN(n662) );
  XNOR2_X1 U745 ( .A(G288), .B(G299), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U747 ( .A(n663), .B(G290), .Z(n664) );
  XNOR2_X1 U748 ( .A(G305), .B(n664), .ZN(n665) );
  XNOR2_X1 U749 ( .A(G166), .B(n665), .ZN(n860) );
  XOR2_X1 U750 ( .A(n860), .B(n666), .Z(n667) );
  NOR2_X1 U751 ( .A1(n669), .A2(n667), .ZN(n671) );
  AND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(KEYINPUT85), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT20), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G235), .A2(G236), .ZN(n677) );
  XOR2_X1 U762 ( .A(KEYINPUT86), .B(n677), .Z(n678) );
  NOR2_X1 U763 ( .A1(G238), .A2(n678), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G57), .A2(n679), .ZN(n838) );
  NAND2_X1 U765 ( .A1(G567), .A2(n838), .ZN(n680) );
  XOR2_X1 U766 ( .A(KEYINPUT87), .B(n680), .Z(n685) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U769 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U770 ( .A1(G96), .A2(n683), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n839), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n906) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n686) );
  XNOR2_X1 U774 ( .A(KEYINPUT88), .B(n686), .ZN(n687) );
  NOR2_X1 U775 ( .A1(n906), .A2(n687), .ZN(n688) );
  XOR2_X1 U776 ( .A(KEYINPUT89), .B(n688), .Z(n837) );
  NAND2_X1 U777 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U778 ( .A1(G102), .A2(n888), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G138), .A2(n889), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U781 ( .A1(G114), .A2(n892), .ZN(n692) );
  NAND2_X1 U782 ( .A1(G126), .A2(n893), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U784 ( .A1(n694), .A2(n693), .ZN(G164) );
  INV_X1 U785 ( .A(G301), .ZN(G171) );
  NAND2_X1 U786 ( .A1(G160), .A2(G40), .ZN(n800) );
  NAND2_X1 U787 ( .A1(KEYINPUT97), .A2(n800), .ZN(n698) );
  INV_X1 U788 ( .A(KEYINPUT97), .ZN(n696) );
  INV_X1 U789 ( .A(n800), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n801) );
  NAND2_X1 U793 ( .A1(G8), .A2(n710), .ZN(n774) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U795 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U796 ( .A1(n774), .A2(n701), .ZN(n779) );
  INV_X1 U797 ( .A(n744), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n702), .A2(G1961), .ZN(n703) );
  XOR2_X1 U799 ( .A(KEYINPUT98), .B(n703), .Z(n705) );
  XNOR2_X1 U800 ( .A(KEYINPUT99), .B(n710), .ZN(n716) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U802 ( .A1(n716), .A2(n946), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n736), .A2(G171), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n716), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U806 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  INV_X1 U807 ( .A(G1956), .ZN(n994) );
  NOR2_X1 U808 ( .A1(n994), .A2(n716), .ZN(n707) );
  NOR2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n725) );
  NOR2_X1 U810 ( .A1(n967), .A2(n725), .ZN(n709) );
  XOR2_X1 U811 ( .A(n709), .B(KEYINPUT28), .Z(n729) );
  INV_X1 U812 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U813 ( .A1(n710), .A2(n942), .ZN(n712) );
  XNOR2_X1 U814 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U815 ( .A1(n744), .A2(G1341), .ZN(n713) );
  NAND2_X1 U816 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U817 ( .A1(n974), .A2(n715), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n722), .A2(n861), .ZN(n720) );
  NAND2_X1 U819 ( .A1(n716), .A2(G2067), .ZN(n718) );
  NAND2_X1 U820 ( .A1(G1348), .A2(n744), .ZN(n717) );
  NAND2_X1 U821 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U822 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U823 ( .A(n721), .B(KEYINPUT100), .ZN(n724) );
  OR2_X1 U824 ( .A1(n722), .A2(n861), .ZN(n723) );
  NAND2_X1 U825 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U826 ( .A1(n967), .A2(n725), .ZN(n726) );
  NAND2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U828 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U829 ( .A(KEYINPUT29), .B(n730), .Z(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n743) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n744), .ZN(n753) );
  NOR2_X1 U832 ( .A1(n756), .A2(n753), .ZN(n733) );
  NAND2_X1 U833 ( .A1(G8), .A2(n521), .ZN(n734) );
  XNOR2_X1 U834 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U835 ( .A1(G168), .A2(n735), .ZN(n738) );
  NOR2_X1 U836 ( .A1(G171), .A2(n736), .ZN(n737) );
  NAND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n754), .A2(G286), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n744), .ZN(n746) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n774), .ZN(n745) );
  NOR2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U842 ( .A1(n747), .A2(G303), .ZN(n748) );
  XOR2_X1 U843 ( .A(KEYINPUT103), .B(n748), .Z(n749) );
  NAND2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n751), .A2(G8), .ZN(n752) );
  XNOR2_X1 U846 ( .A(n752), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(n753), .ZN(n758) );
  INV_X1 U848 ( .A(n754), .ZN(n755) );
  NOR2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n772) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n966), .A2(n761), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n772), .A2(n762), .ZN(n764) );
  NOR2_X1 U856 ( .A1(n774), .A2(n522), .ZN(n763) );
  NOR2_X1 U857 ( .A1(n765), .A2(KEYINPUT33), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n966), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U859 ( .A1(n766), .A2(n774), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U862 ( .A1(n769), .A2(n983), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(n773), .B(KEYINPUT104), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n816) );
  NAND2_X1 U870 ( .A1(n893), .A2(G119), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT91), .B(n780), .Z(n782) );
  NAND2_X1 U872 ( .A1(n892), .A2(G107), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT92), .B(n783), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G95), .A2(n888), .ZN(n785) );
  NAND2_X1 U876 ( .A1(G131), .A2(n889), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n899) );
  XNOR2_X1 U879 ( .A(KEYINPUT93), .B(G1991), .ZN(n947) );
  NOR2_X1 U880 ( .A1(n899), .A2(n947), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G105), .A2(n888), .ZN(n788) );
  XNOR2_X1 U882 ( .A(n788), .B(KEYINPUT38), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G117), .A2(n892), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G129), .A2(n893), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U886 ( .A(KEYINPUT94), .B(n791), .Z(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G141), .A2(n889), .ZN(n794) );
  XNOR2_X1 U889 ( .A(KEYINPUT95), .B(n794), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U891 ( .A(KEYINPUT96), .B(n797), .Z(n881) );
  AND2_X1 U892 ( .A1(G1996), .A2(n881), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n921) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n827) );
  INV_X1 U895 ( .A(n827), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n921), .A2(n802), .ZN(n820) );
  INV_X1 U897 ( .A(n820), .ZN(n813) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n817) );
  NAND2_X1 U899 ( .A1(n889), .A2(G140), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT90), .ZN(n805) );
  NAND2_X1 U901 ( .A1(G104), .A2(n888), .ZN(n804) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U903 ( .A(KEYINPUT34), .B(n806), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G116), .A2(n892), .ZN(n808) );
  NAND2_X1 U905 ( .A1(G128), .A2(n893), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U907 ( .A(KEYINPUT35), .B(n809), .Z(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n812), .ZN(n885) );
  NOR2_X1 U910 ( .A1(n817), .A2(n885), .ZN(n919) );
  NAND2_X1 U911 ( .A1(n827), .A2(n919), .ZN(n825) );
  NAND2_X1 U912 ( .A1(n813), .A2(n825), .ZN(n814) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n965) );
  OR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n817), .A2(n885), .ZN(n920) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n823) );
  AND2_X1 U917 ( .A1(n947), .A2(n899), .ZN(n926) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U919 ( .A1(n926), .A2(n818), .ZN(n819) );
  NOR2_X1 U920 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U921 ( .A1(n881), .A2(G1996), .ZN(n932) );
  NOR2_X1 U922 ( .A1(n821), .A2(n932), .ZN(n822) );
  XOR2_X1 U923 ( .A(n823), .B(n822), .Z(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n920), .A2(n826), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U928 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n832), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n834) );
  INV_X1 U931 ( .A(G661), .ZN(n833) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n835), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U935 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT109), .B(G2090), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n842), .B(G2096), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(G2678), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2100), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U950 ( .A(G2474), .B(G1956), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n851), .B(KEYINPUT110), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U956 ( .A(G1976), .B(G1981), .Z(n855) );
  XNOR2_X1 U957 ( .A(G1961), .B(G1971), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U959 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U960 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(G229) );
  XOR2_X1 U962 ( .A(n860), .B(G286), .Z(n863) );
  XNOR2_X1 U963 ( .A(G301), .B(n861), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n864), .B(n974), .Z(n865) );
  NOR2_X1 U966 ( .A1(G37), .A2(n865), .ZN(G397) );
  NAND2_X1 U967 ( .A1(G100), .A2(n888), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G112), .A2(n892), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT112), .B(n868), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n893), .A2(G124), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G136), .A2(n889), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G118), .A2(n892), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G130), .A2(n893), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n888), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G142), .A2(n889), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n884) );
  XNOR2_X1 U984 ( .A(G160), .B(n881), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n882), .B(G162), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n885), .B(n927), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n904) );
  XOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n901) );
  NAND2_X1 U990 ( .A1(G103), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G115), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G127), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n914) );
  XNOR2_X1 U998 ( .A(n899), .B(n914), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(G164), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT108), .B(n906), .Z(G319) );
  XNOR2_X1 U1004 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(KEYINPUT114), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n913), .A2(G319), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1014 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1025) );
  INV_X1 U1015 ( .A(KEYINPUT55), .ZN(n939) );
  XOR2_X1 U1016 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n937) );
  XOR2_X1 U1017 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n917), .Z(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n923) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT115), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n937), .B(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(G2090), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(G35), .ZN(n960) );
  XNOR2_X1 U1038 ( .A(G32), .B(n942), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n951) );
  XOR2_X1 U1043 ( .A(n946), .B(G27), .Z(n949) );
  XOR2_X1 U1044 ( .A(n947), .B(G25), .Z(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n954), .B(KEYINPUT53), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(n955), .B(KEYINPUT118), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G2084), .B(G34), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT55), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n963), .B(KEYINPUT119), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n964), .ZN(n1021) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  NOR2_X1 U1059 ( .A1(n522), .A2(n965), .ZN(n973) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT123), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n967), .B(G1956), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G303), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n974), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n989) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1348), .B(KEYINPUT121), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(KEYINPUT122), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n982), .B(KEYINPUT120), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n1019) );
  INV_X1 U1080 ( .A(G16), .ZN(n1017) );
  XOR2_X1 U1081 ( .A(G4), .B(KEYINPUT124), .Z(n993) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n993), .B(n992), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G20), .B(n994), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT125), .B(n1001), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1002), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G5), .B(G1961), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G1986), .B(KEYINPUT126), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(G24), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1025), .B(n1024), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

